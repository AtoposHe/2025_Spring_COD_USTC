
`timescale 1ns/1ps
module mem_bram #(
    parameter ADDR_WIDTH = 10,		//地址宽度
    parameter DATA_WIDTH = 128		//数据宽度
)(
    input                   clk,   // Clock
    input [ADDR_WIDTH-1:0]  raddr,  // Address
    input [ADDR_WIDTH-1:0]  waddr,  // Address
    input [DATA_WIDTH-1:0]  din,   // Data Input
    input                   we,    // Write Enable
    output [DATA_WIDTH-1:0] dout   // Data Output
); 
    reg [ADDR_WIDTH-1:0] addr_r;  // Address Register
    reg [DATA_WIDTH-1:0] ram [0:(1 << ADDR_WIDTH)-1];
    integer i;
    initial begin
        ram[0][31:0] = 32'd1052567479;
        ram[0][63:32] = 32'd3962591981;
        ram[0][95:64] = 32'd3364158968;
        ram[0][127:96] = 32'd2890460227;
        ram[1][31:0] = 32'd3294865998;
        ram[1][63:32] = 32'd3904772148;
        ram[1][95:64] = 32'd4003091934;
        ram[1][127:96] = 32'd3045195451;
        ram[2][31:0] = 32'd606447009;
        ram[2][63:32] = 32'd1508884471;
        ram[2][95:64] = 32'd2855376560;
        ram[2][127:96] = 32'd2135414422;
        ram[3][31:0] = 32'd770777372;
        ram[3][63:32] = 32'd675467997;
        ram[3][95:64] = 32'd1785532064;
        ram[3][127:96] = 32'd440331261;
        ram[4][31:0] = 32'd1426394555;
        ram[4][63:32] = 32'd713149634;
        ram[4][95:64] = 32'd3721935424;
        ram[4][127:96] = 32'd694124835;
        ram[5][31:0] = 32'd3887719615;
        ram[5][63:32] = 32'd2131512427;
        ram[5][95:64] = 32'd3582627947;
        ram[5][127:96] = 32'd789024827;
        ram[6][31:0] = 32'd1235305684;
        ram[6][63:32] = 32'd3096215726;
        ram[6][95:64] = 32'd59093393;
        ram[6][127:96] = 32'd1793516677;
        ram[7][31:0] = 32'd3711284261;
        ram[7][63:32] = 32'd233984458;
        ram[7][95:64] = 32'd280682631;
        ram[7][127:96] = 32'd3024886858;
        ram[8][31:0] = 32'd3943143764;
        ram[8][63:32] = 32'd437396483;
        ram[8][95:64] = 32'd3140383792;
        ram[8][127:96] = 32'd3596422925;
        ram[9][31:0] = 32'd3203529788;
        ram[9][63:32] = 32'd1883382384;
        ram[9][95:64] = 32'd1832735743;
        ram[9][127:96] = 32'd2778868458;
        ram[10][31:0] = 32'd334310572;
        ram[10][63:32] = 32'd547420335;
        ram[10][95:64] = 32'd631245937;
        ram[10][127:96] = 32'd2262236211;
        ram[11][31:0] = 32'd2295093428;
        ram[11][63:32] = 32'd3807651913;
        ram[11][95:64] = 32'd3718565962;
        ram[11][127:96] = 32'd456343954;
        ram[12][31:0] = 32'd3884411445;
        ram[12][63:32] = 32'd4260315682;
        ram[12][95:64] = 32'd317339329;
        ram[12][127:96] = 32'd2846119786;
        ram[13][31:0] = 32'd2810219511;
        ram[13][63:32] = 32'd4067531662;
        ram[13][95:64] = 32'd1273374471;
        ram[13][127:96] = 32'd855085249;
        ram[14][31:0] = 32'd2040694399;
        ram[14][63:32] = 32'd3664626015;
        ram[14][95:64] = 32'd1265219196;
        ram[14][127:96] = 32'd482179054;
        ram[15][31:0] = 32'd1557958011;
        ram[15][63:32] = 32'd468031354;
        ram[15][95:64] = 32'd317058348;
        ram[15][127:96] = 32'd812315635;
        ram[16][31:0] = 32'd819283579;
        ram[16][63:32] = 32'd1536885837;
        ram[16][95:64] = 32'd2714239827;
        ram[16][127:96] = 32'd3494148640;
        ram[17][31:0] = 32'd88490023;
        ram[17][63:32] = 32'd2018933038;
        ram[17][95:64] = 32'd1396858963;
        ram[17][127:96] = 32'd3173125001;
        ram[18][31:0] = 32'd1361381559;
        ram[18][63:32] = 32'd546788671;
        ram[18][95:64] = 32'd2836015271;
        ram[18][127:96] = 32'd1791303464;
        ram[19][31:0] = 32'd3925384761;
        ram[19][63:32] = 32'd3109637631;
        ram[19][95:64] = 32'd728046435;
        ram[19][127:96] = 32'd3294863484;
        ram[20][31:0] = 32'd1142305230;
        ram[20][63:32] = 32'd1252273539;
        ram[20][95:64] = 32'd1161768830;
        ram[20][127:96] = 32'd4103514108;
        ram[21][31:0] = 32'd3678239471;
        ram[21][63:32] = 32'd3558159285;
        ram[21][95:64] = 32'd2026415795;
        ram[21][127:96] = 32'd2832515348;
        ram[22][31:0] = 32'd4180574515;
        ram[22][63:32] = 32'd777576892;
        ram[22][95:64] = 32'd610397100;
        ram[22][127:96] = 32'd1707606940;
        ram[23][31:0] = 32'd732174983;
        ram[23][63:32] = 32'd3982696287;
        ram[23][95:64] = 32'd4279075714;
        ram[23][127:96] = 32'd4186162648;
        ram[24][31:0] = 32'd3668307642;
        ram[24][63:32] = 32'd1844783002;
        ram[24][95:64] = 32'd2262198691;
        ram[24][127:96] = 32'd1962326579;
        ram[25][31:0] = 32'd2509988248;
        ram[25][63:32] = 32'd3945960348;
        ram[25][95:64] = 32'd2639049148;
        ram[25][127:96] = 32'd1753914851;
        ram[26][31:0] = 32'd2137822137;
        ram[26][63:32] = 32'd2079086660;
        ram[26][95:64] = 32'd1346540745;
        ram[26][127:96] = 32'd2778245487;
        ram[27][31:0] = 32'd3644488255;
        ram[27][63:32] = 32'd664815512;
        ram[27][95:64] = 32'd3750726883;
        ram[27][127:96] = 32'd2870920926;
        ram[28][31:0] = 32'd53516149;
        ram[28][63:32] = 32'd2628436063;
        ram[28][95:64] = 32'd574419132;
        ram[28][127:96] = 32'd1787837868;
        ram[29][31:0] = 32'd232587118;
        ram[29][63:32] = 32'd222685664;
        ram[29][95:64] = 32'd3910724969;
        ram[29][127:96] = 32'd2347492591;
        ram[30][31:0] = 32'd3159296284;
        ram[30][63:32] = 32'd1116625760;
        ram[30][95:64] = 32'd2382385405;
        ram[30][127:96] = 32'd2378157637;
        ram[31][31:0] = 32'd695025908;
        ram[31][63:32] = 32'd1547082423;
        ram[31][95:64] = 32'd2166982801;
        ram[31][127:96] = 32'd1861995505;
        ram[32][31:0] = 32'd2999443473;
        ram[32][63:32] = 32'd4213028843;
        ram[32][95:64] = 32'd1440556275;
        ram[32][127:96] = 32'd3900854079;
        ram[33][31:0] = 32'd1523580593;
        ram[33][63:32] = 32'd2214113554;
        ram[33][95:64] = 32'd137763915;
        ram[33][127:96] = 32'd1164078325;
        ram[34][31:0] = 32'd796988188;
        ram[34][63:32] = 32'd2021339031;
        ram[34][95:64] = 32'd2736216411;
        ram[34][127:96] = 32'd932387086;
        ram[35][31:0] = 32'd3627393903;
        ram[35][63:32] = 32'd1824634388;
        ram[35][95:64] = 32'd662381207;
        ram[35][127:96] = 32'd3652162657;
        ram[36][31:0] = 32'd3389748868;
        ram[36][63:32] = 32'd3995848082;
        ram[36][95:64] = 32'd1744338134;
        ram[36][127:96] = 32'd3842886285;
        ram[37][31:0] = 32'd1157076026;
        ram[37][63:32] = 32'd3091660807;
        ram[37][95:64] = 32'd2857650347;
        ram[37][127:96] = 32'd1274566182;
        ram[38][31:0] = 32'd1978607299;
        ram[38][63:32] = 32'd3554490906;
        ram[38][95:64] = 32'd3756857754;
        ram[38][127:96] = 32'd2556299901;
        ram[39][31:0] = 32'd3397644777;
        ram[39][63:32] = 32'd295494249;
        ram[39][95:64] = 32'd3357021415;
        ram[39][127:96] = 32'd885040515;
        ram[40][31:0] = 32'd688845184;
        ram[40][63:32] = 32'd1723706081;
        ram[40][95:64] = 32'd262508675;
        ram[40][127:96] = 32'd120689546;
        ram[41][31:0] = 32'd10763549;
        ram[41][63:32] = 32'd3249592251;
        ram[41][95:64] = 32'd1582126961;
        ram[41][127:96] = 32'd3262096531;
        ram[42][31:0] = 32'd3104257694;
        ram[42][63:32] = 32'd1157869169;
        ram[42][95:64] = 32'd4056548843;
        ram[42][127:96] = 32'd516640682;
        ram[43][31:0] = 32'd909425390;
        ram[43][63:32] = 32'd3560746765;
        ram[43][95:64] = 32'd2494804107;
        ram[43][127:96] = 32'd1660422906;
        ram[44][31:0] = 32'd1240149642;
        ram[44][63:32] = 32'd1530014160;
        ram[44][95:64] = 32'd2218298793;
        ram[44][127:96] = 32'd2165023982;
        ram[45][31:0] = 32'd1394926462;
        ram[45][63:32] = 32'd1038253186;
        ram[45][95:64] = 32'd830768617;
        ram[45][127:96] = 32'd309566207;
        ram[46][31:0] = 32'd2586566993;
        ram[46][63:32] = 32'd4181767754;
        ram[46][95:64] = 32'd3269096103;
        ram[46][127:96] = 32'd579136898;
        ram[47][31:0] = 32'd3715826206;
        ram[47][63:32] = 32'd1457465443;
        ram[47][95:64] = 32'd1159409871;
        ram[47][127:96] = 32'd3285354185;
        ram[48][31:0] = 32'd251807735;
        ram[48][63:32] = 32'd389818431;
        ram[48][95:64] = 32'd1081961558;
        ram[48][127:96] = 32'd1068866777;
        ram[49][31:0] = 32'd871728998;
        ram[49][63:32] = 32'd3233146207;
        ram[49][95:64] = 32'd1825329058;
        ram[49][127:96] = 32'd80750494;
        ram[50][31:0] = 32'd2827824628;
        ram[50][63:32] = 32'd1105729140;
        ram[50][95:64] = 32'd1009518837;
        ram[50][127:96] = 32'd1252458418;
        ram[51][31:0] = 32'd1243827460;
        ram[51][63:32] = 32'd2438118847;
        ram[51][95:64] = 32'd617153583;
        ram[51][127:96] = 32'd867306624;
        ram[52][31:0] = 32'd1518584672;
        ram[52][63:32] = 32'd2811362265;
        ram[52][95:64] = 32'd1216497215;
        ram[52][127:96] = 32'd2113102357;
        ram[53][31:0] = 32'd3427452440;
        ram[53][63:32] = 32'd3842928591;
        ram[53][95:64] = 32'd67071196;
        ram[53][127:96] = 32'd1968456532;
        ram[54][31:0] = 32'd3763448983;
        ram[54][63:32] = 32'd91812431;
        ram[54][95:64] = 32'd709857341;
        ram[54][127:96] = 32'd2119043502;
        ram[55][31:0] = 32'd3956104701;
        ram[55][63:32] = 32'd3402247746;
        ram[55][95:64] = 32'd128119112;
        ram[55][127:96] = 32'd1645865683;
        ram[56][31:0] = 32'd1160411914;
        ram[56][63:32] = 32'd638184484;
        ram[56][95:64] = 32'd2785708549;
        ram[56][127:96] = 32'd3087655498;
        ram[57][31:0] = 32'd1874932830;
        ram[57][63:32] = 32'd3060630889;
        ram[57][95:64] = 32'd377097911;
        ram[57][127:96] = 32'd528724415;
        ram[58][31:0] = 32'd4268345978;
        ram[58][63:32] = 32'd4110817650;
        ram[58][95:64] = 32'd1388060105;
        ram[58][127:96] = 32'd483824422;
        ram[59][31:0] = 32'd2037725383;
        ram[59][63:32] = 32'd1838823857;
        ram[59][95:64] = 32'd3263906087;
        ram[59][127:96] = 32'd777675197;
        ram[60][31:0] = 32'd2405468028;
        ram[60][63:32] = 32'd2418047968;
        ram[60][95:64] = 32'd1678087538;
        ram[60][127:96] = 32'd975543220;
        ram[61][31:0] = 32'd1765401337;
        ram[61][63:32] = 32'd1169530796;
        ram[61][95:64] = 32'd2920595436;
        ram[61][127:96] = 32'd3098617292;
        ram[62][31:0] = 32'd567480644;
        ram[62][63:32] = 32'd1695986456;
        ram[62][95:64] = 32'd1214633845;
        ram[62][127:96] = 32'd2582319262;
        ram[63][31:0] = 32'd1646463308;
        ram[63][63:32] = 32'd3083274420;
        ram[63][95:64] = 32'd2992602956;
        ram[63][127:96] = 32'd3333567760;
        ram[64][31:0] = 32'd2873197191;
        ram[64][63:32] = 32'd1521182444;
        ram[64][95:64] = 32'd2245328102;
        ram[64][127:96] = 32'd964259512;
        ram[65][31:0] = 32'd3678551605;
        ram[65][63:32] = 32'd1946819819;
        ram[65][95:64] = 32'd1949534506;
        ram[65][127:96] = 32'd1923525205;
        ram[66][31:0] = 32'd3744119204;
        ram[66][63:32] = 32'd4016900671;
        ram[66][95:64] = 32'd1955864689;
        ram[66][127:96] = 32'd2586515488;
        ram[67][31:0] = 32'd1722456956;
        ram[67][63:32] = 32'd221469839;
        ram[67][95:64] = 32'd3591863440;
        ram[67][127:96] = 32'd4184036158;
        ram[68][31:0] = 32'd2613524396;
        ram[68][63:32] = 32'd262445657;
        ram[68][95:64] = 32'd1993005996;
        ram[68][127:96] = 32'd1691264788;
        ram[69][31:0] = 32'd1830683552;
        ram[69][63:32] = 32'd2186026964;
        ram[69][95:64] = 32'd2738662472;
        ram[69][127:96] = 32'd1394720320;
        ram[70][31:0] = 32'd778579737;
        ram[70][63:32] = 32'd2713817115;
        ram[70][95:64] = 32'd643220710;
        ram[70][127:96] = 32'd2130912552;
        ram[71][31:0] = 32'd450921526;
        ram[71][63:32] = 32'd2092726877;
        ram[71][95:64] = 32'd782042751;
        ram[71][127:96] = 32'd3656423157;
        ram[72][31:0] = 32'd2987361026;
        ram[72][63:32] = 32'd3503208650;
        ram[72][95:64] = 32'd193368078;
        ram[72][127:96] = 32'd1270361158;
        ram[73][31:0] = 32'd2882588279;
        ram[73][63:32] = 32'd3661832280;
        ram[73][95:64] = 32'd1462825451;
        ram[73][127:96] = 32'd2157362138;
        ram[74][31:0] = 32'd2438739140;
        ram[74][63:32] = 32'd1173911246;
        ram[74][95:64] = 32'd2569764979;
        ram[74][127:96] = 32'd205743923;
        ram[75][31:0] = 32'd3464558724;
        ram[75][63:32] = 32'd3805465914;
        ram[75][95:64] = 32'd1757630826;
        ram[75][127:96] = 32'd756679895;
        ram[76][31:0] = 32'd3131755163;
        ram[76][63:32] = 32'd2985268612;
        ram[76][95:64] = 32'd2048220064;
        ram[76][127:96] = 32'd395268976;
        ram[77][31:0] = 32'd1555365123;
        ram[77][63:32] = 32'd1157989693;
        ram[77][95:64] = 32'd892285550;
        ram[77][127:96] = 32'd757719279;
        ram[78][31:0] = 32'd2911720261;
        ram[78][63:32] = 32'd2709848361;
        ram[78][95:64] = 32'd672074592;
        ram[78][127:96] = 32'd1958764270;
        ram[79][31:0] = 32'd2469986364;
        ram[79][63:32] = 32'd1975671844;
        ram[79][95:64] = 32'd3064576727;
        ram[79][127:96] = 32'd3883511213;
        ram[80][31:0] = 32'd2659365932;
        ram[80][63:32] = 32'd2227829365;
        ram[80][95:64] = 32'd1384846976;
        ram[80][127:96] = 32'd200882046;
        ram[81][31:0] = 32'd2565321190;
        ram[81][63:32] = 32'd2573803079;
        ram[81][95:64] = 32'd4237884957;
        ram[81][127:96] = 32'd192410890;
        ram[82][31:0] = 32'd3264070670;
        ram[82][63:32] = 32'd3283575319;
        ram[82][95:64] = 32'd19614130;
        ram[82][127:96] = 32'd2981950880;
        ram[83][31:0] = 32'd4118120138;
        ram[83][63:32] = 32'd3504452332;
        ram[83][95:64] = 32'd1684630731;
        ram[83][127:96] = 32'd459514534;
        ram[84][31:0] = 32'd966779298;
        ram[84][63:32] = 32'd4218420959;
        ram[84][95:64] = 32'd2832891657;
        ram[84][127:96] = 32'd3901609669;
        ram[85][31:0] = 32'd2309224711;
        ram[85][63:32] = 32'd1297508340;
        ram[85][95:64] = 32'd3867550255;
        ram[85][127:96] = 32'd4268882280;
        ram[86][31:0] = 32'd100362266;
        ram[86][63:32] = 32'd2316252777;
        ram[86][95:64] = 32'd2418381156;
        ram[86][127:96] = 32'd3975745931;
        ram[87][31:0] = 32'd2859983252;
        ram[87][63:32] = 32'd2089693596;
        ram[87][95:64] = 32'd1993790010;
        ram[87][127:96] = 32'd1483615543;
        ram[88][31:0] = 32'd2089405516;
        ram[88][63:32] = 32'd1007787516;
        ram[88][95:64] = 32'd4104199402;
        ram[88][127:96] = 32'd4231388117;
        ram[89][31:0] = 32'd328648182;
        ram[89][63:32] = 32'd2244387970;
        ram[89][95:64] = 32'd2281669903;
        ram[89][127:96] = 32'd3857920595;
        ram[90][31:0] = 32'd1685941148;
        ram[90][63:32] = 32'd3332500024;
        ram[90][95:64] = 32'd2761902832;
        ram[90][127:96] = 32'd803716268;
        ram[91][31:0] = 32'd3270560608;
        ram[91][63:32] = 32'd92649394;
        ram[91][95:64] = 32'd4105913331;
        ram[91][127:96] = 32'd3378755930;
        ram[92][31:0] = 32'd3625661537;
        ram[92][63:32] = 32'd2921962052;
        ram[92][95:64] = 32'd1101997953;
        ram[92][127:96] = 32'd3980939607;
        ram[93][31:0] = 32'd1069657798;
        ram[93][63:32] = 32'd2879679012;
        ram[93][95:64] = 32'd276518235;
        ram[93][127:96] = 32'd86563587;
        ram[94][31:0] = 32'd2007598323;
        ram[94][63:32] = 32'd2225356755;
        ram[94][95:64] = 32'd1683535556;
        ram[94][127:96] = 32'd203189148;
        ram[95][31:0] = 32'd2016133482;
        ram[95][63:32] = 32'd1644109573;
        ram[95][95:64] = 32'd246575701;
        ram[95][127:96] = 32'd1470696070;
        ram[96][31:0] = 32'd1338121990;
        ram[96][63:32] = 32'd1312176869;
        ram[96][95:64] = 32'd3060009435;
        ram[96][127:96] = 32'd1682531476;
        ram[97][31:0] = 32'd3061490345;
        ram[97][63:32] = 32'd3581898418;
        ram[97][95:64] = 32'd2619734395;
        ram[97][127:96] = 32'd215431964;
        ram[98][31:0] = 32'd4014398129;
        ram[98][63:32] = 32'd1253624254;
        ram[98][95:64] = 32'd3249060309;
        ram[98][127:96] = 32'd960981275;
        ram[99][31:0] = 32'd1974444420;
        ram[99][63:32] = 32'd2655648054;
        ram[99][95:64] = 32'd3583158237;
        ram[99][127:96] = 32'd1694067374;
        ram[100][31:0] = 32'd2624678043;
        ram[100][63:32] = 32'd1181135291;
        ram[100][95:64] = 32'd1240298673;
        ram[100][127:96] = 32'd1230970457;
        ram[101][31:0] = 32'd2974441075;
        ram[101][63:32] = 32'd1501224403;
        ram[101][95:64] = 32'd3598914984;
        ram[101][127:96] = 32'd2926448752;
        ram[102][31:0] = 32'd2708666325;
        ram[102][63:32] = 32'd664332654;
        ram[102][95:64] = 32'd2554823396;
        ram[102][127:96] = 32'd1912192808;
        ram[103][31:0] = 32'd251190816;
        ram[103][63:32] = 32'd42785687;
        ram[103][95:64] = 32'd791976254;
        ram[103][127:96] = 32'd3418827215;
        ram[104][31:0] = 32'd3371794246;
        ram[104][63:32] = 32'd3457950605;
        ram[104][95:64] = 32'd3358504200;
        ram[104][127:96] = 32'd3137721503;
        ram[105][31:0] = 32'd3236855211;
        ram[105][63:32] = 32'd3199121285;
        ram[105][95:64] = 32'd4144966284;
        ram[105][127:96] = 32'd2356837183;
        ram[106][31:0] = 32'd2630810105;
        ram[106][63:32] = 32'd2959861491;
        ram[106][95:64] = 32'd4113724443;
        ram[106][127:96] = 32'd3990194643;
        ram[107][31:0] = 32'd3112127436;
        ram[107][63:32] = 32'd3410880727;
        ram[107][95:64] = 32'd3912201120;
        ram[107][127:96] = 32'd1792006120;
        ram[108][31:0] = 32'd807161466;
        ram[108][63:32] = 32'd363795349;
        ram[108][95:64] = 32'd1755049189;
        ram[108][127:96] = 32'd2035856504;
        ram[109][31:0] = 32'd2811885061;
        ram[109][63:32] = 32'd1332405155;
        ram[109][95:64] = 32'd873569353;
        ram[109][127:96] = 32'd1956260871;
        ram[110][31:0] = 32'd2562872072;
        ram[110][63:32] = 32'd65904936;
        ram[110][95:64] = 32'd1741314760;
        ram[110][127:96] = 32'd3927924680;
        ram[111][31:0] = 32'd4084632541;
        ram[111][63:32] = 32'd3196251038;
        ram[111][95:64] = 32'd3408163439;
        ram[111][127:96] = 32'd1208282183;
        ram[112][31:0] = 32'd1265298441;
        ram[112][63:32] = 32'd2908833870;
        ram[112][95:64] = 32'd2162667854;
        ram[112][127:96] = 32'd1966989712;
        ram[113][31:0] = 32'd660059285;
        ram[113][63:32] = 32'd285543293;
        ram[113][95:64] = 32'd2191347482;
        ram[113][127:96] = 32'd2580577157;
        ram[114][31:0] = 32'd321448812;
        ram[114][63:32] = 32'd2500934454;
        ram[114][95:64] = 32'd2264632454;
        ram[114][127:96] = 32'd1531900981;
        ram[115][31:0] = 32'd2220856156;
        ram[115][63:32] = 32'd3428994727;
        ram[115][95:64] = 32'd1385003637;
        ram[115][127:96] = 32'd4166078644;
        ram[116][31:0] = 32'd1092151286;
        ram[116][63:32] = 32'd3508624685;
        ram[116][95:64] = 32'd3264154007;
        ram[116][127:96] = 32'd1066574642;
        ram[117][31:0] = 32'd1244655582;
        ram[117][63:32] = 32'd4275884649;
        ram[117][95:64] = 32'd1434334882;
        ram[117][127:96] = 32'd3824336063;
        ram[118][31:0] = 32'd4261511285;
        ram[118][63:32] = 32'd3858581669;
        ram[118][95:64] = 32'd1723651348;
        ram[118][127:96] = 32'd3328634438;
        ram[119][31:0] = 32'd2866816344;
        ram[119][63:32] = 32'd3782855187;
        ram[119][95:64] = 32'd1734380702;
        ram[119][127:96] = 32'd4019054393;
        ram[120][31:0] = 32'd799026300;
        ram[120][63:32] = 32'd3611509395;
        ram[120][95:64] = 32'd2956058280;
        ram[120][127:96] = 32'd3314459181;
        ram[121][31:0] = 32'd1119167468;
        ram[121][63:32] = 32'd453359906;
        ram[121][95:64] = 32'd3122163460;
        ram[121][127:96] = 32'd53661114;
        ram[122][31:0] = 32'd1111823230;
        ram[122][63:32] = 32'd1327010194;
        ram[122][95:64] = 32'd1847146603;
        ram[122][127:96] = 32'd2232007344;
        ram[123][31:0] = 32'd2825740953;
        ram[123][63:32] = 32'd3318295190;
        ram[123][95:64] = 32'd2219142457;
        ram[123][127:96] = 32'd2985661865;
        ram[124][31:0] = 32'd3672699243;
        ram[124][63:32] = 32'd253968604;
        ram[124][95:64] = 32'd920808543;
        ram[124][127:96] = 32'd3119393922;
        ram[125][31:0] = 32'd705804285;
        ram[125][63:32] = 32'd4273805406;
        ram[125][95:64] = 32'd2172460038;
        ram[125][127:96] = 32'd2038481495;
        ram[126][31:0] = 32'd1574083226;
        ram[126][63:32] = 32'd3731120467;
        ram[126][95:64] = 32'd799205872;
        ram[126][127:96] = 32'd3526605853;
        ram[127][31:0] = 32'd3420814826;
        ram[127][63:32] = 32'd282828349;
        ram[127][95:64] = 32'd636963736;
        ram[127][127:96] = 32'd667745192;
        ram[128][31:0] = 32'd3815785216;
        ram[128][63:32] = 32'd444266860;
        ram[128][95:64] = 32'd3329925324;
        ram[128][127:96] = 32'd2421804531;
        ram[129][31:0] = 32'd44690167;
        ram[129][63:32] = 32'd4145418118;
        ram[129][95:64] = 32'd1018664874;
        ram[129][127:96] = 32'd1574109177;
        ram[130][31:0] = 32'd847712690;
        ram[130][63:32] = 32'd3118728776;
        ram[130][95:64] = 32'd684068191;
        ram[130][127:96] = 32'd40985424;
        ram[131][31:0] = 32'd3607396520;
        ram[131][63:32] = 32'd3236712843;
        ram[131][95:64] = 32'd3914327828;
        ram[131][127:96] = 32'd66118690;
        ram[132][31:0] = 32'd4235592281;
        ram[132][63:32] = 32'd1798434561;
        ram[132][95:64] = 32'd197641397;
        ram[132][127:96] = 32'd1917508662;
        ram[133][31:0] = 32'd2986500363;
        ram[133][63:32] = 32'd998652042;
        ram[133][95:64] = 32'd1477567924;
        ram[133][127:96] = 32'd740792702;
        ram[134][31:0] = 32'd1359838887;
        ram[134][63:32] = 32'd1119348756;
        ram[134][95:64] = 32'd3271843031;
        ram[134][127:96] = 32'd276712892;
        ram[135][31:0] = 32'd3375317644;
        ram[135][63:32] = 32'd239769310;
        ram[135][95:64] = 32'd142287012;
        ram[135][127:96] = 32'd4225807241;
        ram[136][31:0] = 32'd3366506315;
        ram[136][63:32] = 32'd2345963143;
        ram[136][95:64] = 32'd3228427618;
        ram[136][127:96] = 32'd163397476;
        ram[137][31:0] = 32'd1948542852;
        ram[137][63:32] = 32'd4281859846;
        ram[137][95:64] = 32'd3804497467;
        ram[137][127:96] = 32'd2242960485;
        ram[138][31:0] = 32'd822192939;
        ram[138][63:32] = 32'd816505272;
        ram[138][95:64] = 32'd279679526;
        ram[138][127:96] = 32'd3894035056;
        ram[139][31:0] = 32'd2385157507;
        ram[139][63:32] = 32'd3787715714;
        ram[139][95:64] = 32'd762053316;
        ram[139][127:96] = 32'd3250198723;
        ram[140][31:0] = 32'd3966735267;
        ram[140][63:32] = 32'd720640157;
        ram[140][95:64] = 32'd3211385674;
        ram[140][127:96] = 32'd2283251439;
        ram[141][31:0] = 32'd589376832;
        ram[141][63:32] = 32'd1424860412;
        ram[141][95:64] = 32'd4203930147;
        ram[141][127:96] = 32'd3250113416;
        ram[142][31:0] = 32'd74969035;
        ram[142][63:32] = 32'd3416048394;
        ram[142][95:64] = 32'd3977968930;
        ram[142][127:96] = 32'd3866372985;
        ram[143][31:0] = 32'd446317660;
        ram[143][63:32] = 32'd667426504;
        ram[143][95:64] = 32'd277213762;
        ram[143][127:96] = 32'd2498279954;
        ram[144][31:0] = 32'd3483067739;
        ram[144][63:32] = 32'd474077448;
        ram[144][95:64] = 32'd2578797357;
        ram[144][127:96] = 32'd2429845848;
        ram[145][31:0] = 32'd3083515047;
        ram[145][63:32] = 32'd3064431451;
        ram[145][95:64] = 32'd2220997705;
        ram[145][127:96] = 32'd2367557065;
        ram[146][31:0] = 32'd1690895911;
        ram[146][63:32] = 32'd3545634013;
        ram[146][95:64] = 32'd3351735354;
        ram[146][127:96] = 32'd291280601;
        ram[147][31:0] = 32'd228267201;
        ram[147][63:32] = 32'd1882228859;
        ram[147][95:64] = 32'd2568663595;
        ram[147][127:96] = 32'd4103338995;
        ram[148][31:0] = 32'd3890705901;
        ram[148][63:32] = 32'd58166058;
        ram[148][95:64] = 32'd605388411;
        ram[148][127:96] = 32'd4101054525;
        ram[149][31:0] = 32'd3005148523;
        ram[149][63:32] = 32'd3336186297;
        ram[149][95:64] = 32'd901281216;
        ram[149][127:96] = 32'd4293738456;
        ram[150][31:0] = 32'd508264472;
        ram[150][63:32] = 32'd2571072663;
        ram[150][95:64] = 32'd2987575655;
        ram[150][127:96] = 32'd3930150954;
        ram[151][31:0] = 32'd1222723850;
        ram[151][63:32] = 32'd3919297631;
        ram[151][95:64] = 32'd242612497;
        ram[151][127:96] = 32'd172581437;
        ram[152][31:0] = 32'd4136444716;
        ram[152][63:32] = 32'd3925486970;
        ram[152][95:64] = 32'd3603903628;
        ram[152][127:96] = 32'd2389840076;
        ram[153][31:0] = 32'd1075777044;
        ram[153][63:32] = 32'd2147567015;
        ram[153][95:64] = 32'd2943240457;
        ram[153][127:96] = 32'd2283134385;
        ram[154][31:0] = 32'd1433995368;
        ram[154][63:32] = 32'd2569428065;
        ram[154][95:64] = 32'd1302725125;
        ram[154][127:96] = 32'd3667454584;
        ram[155][31:0] = 32'd2816982930;
        ram[155][63:32] = 32'd3470453698;
        ram[155][95:64] = 32'd3878932875;
        ram[155][127:96] = 32'd1284144988;
        ram[156][31:0] = 32'd2824885127;
        ram[156][63:32] = 32'd3903890825;
        ram[156][95:64] = 32'd2443222463;
        ram[156][127:96] = 32'd207512883;
        ram[157][31:0] = 32'd390612325;
        ram[157][63:32] = 32'd3640747;
        ram[157][95:64] = 32'd2440170518;
        ram[157][127:96] = 32'd243801277;
        ram[158][31:0] = 32'd1454516492;
        ram[158][63:32] = 32'd3766781495;
        ram[158][95:64] = 32'd941110408;
        ram[158][127:96] = 32'd2142044604;
        ram[159][31:0] = 32'd3358336986;
        ram[159][63:32] = 32'd2915264513;
        ram[159][95:64] = 32'd2786119313;
        ram[159][127:96] = 32'd343353612;
        ram[160][31:0] = 32'd1294707516;
        ram[160][63:32] = 32'd263459559;
        ram[160][95:64] = 32'd1917049000;
        ram[160][127:96] = 32'd2925530671;
        ram[161][31:0] = 32'd3042117089;
        ram[161][63:32] = 32'd3539970854;
        ram[161][95:64] = 32'd3351083848;
        ram[161][127:96] = 32'd3098822722;
        ram[162][31:0] = 32'd320726234;
        ram[162][63:32] = 32'd2831991724;
        ram[162][95:64] = 32'd3593391115;
        ram[162][127:96] = 32'd2684155943;
        ram[163][31:0] = 32'd441036182;
        ram[163][63:32] = 32'd2986341452;
        ram[163][95:64] = 32'd266085065;
        ram[163][127:96] = 32'd763025037;
        ram[164][31:0] = 32'd3629056107;
        ram[164][63:32] = 32'd668982047;
        ram[164][95:64] = 32'd2565372091;
        ram[164][127:96] = 32'd1343443381;
        ram[165][31:0] = 32'd287497666;
        ram[165][63:32] = 32'd4220104399;
        ram[165][95:64] = 32'd3965663817;
        ram[165][127:96] = 32'd372966818;
        ram[166][31:0] = 32'd1304378213;
        ram[166][63:32] = 32'd2034289997;
        ram[166][95:64] = 32'd4072192775;
        ram[166][127:96] = 32'd2563820725;
        ram[167][31:0] = 32'd3382879701;
        ram[167][63:32] = 32'd3165934849;
        ram[167][95:64] = 32'd2503869172;
        ram[167][127:96] = 32'd222714301;
        ram[168][31:0] = 32'd336862564;
        ram[168][63:32] = 32'd4240157953;
        ram[168][95:64] = 32'd602961986;
        ram[168][127:96] = 32'd953773948;
        ram[169][31:0] = 32'd1873765848;
        ram[169][63:32] = 32'd2364878071;
        ram[169][95:64] = 32'd2364391312;
        ram[169][127:96] = 32'd3630532157;
        ram[170][31:0] = 32'd708134854;
        ram[170][63:32] = 32'd2488012861;
        ram[170][95:64] = 32'd2655148014;
        ram[170][127:96] = 32'd3868012904;
        ram[171][31:0] = 32'd878735113;
        ram[171][63:32] = 32'd1269636871;
        ram[171][95:64] = 32'd3201733946;
        ram[171][127:96] = 32'd1463662090;
        ram[172][31:0] = 32'd2462885890;
        ram[172][63:32] = 32'd743705583;
        ram[172][95:64] = 32'd2378395861;
        ram[172][127:96] = 32'd1508790809;
        ram[173][31:0] = 32'd735552833;
        ram[173][63:32] = 32'd821766607;
        ram[173][95:64] = 32'd3269737490;
        ram[173][127:96] = 32'd688799337;
        ram[174][31:0] = 32'd1822071661;
        ram[174][63:32] = 32'd1856755845;
        ram[174][95:64] = 32'd956868412;
        ram[174][127:96] = 32'd507075352;
        ram[175][31:0] = 32'd1049995550;
        ram[175][63:32] = 32'd2591022462;
        ram[175][95:64] = 32'd2452957524;
        ram[175][127:96] = 32'd2083865596;
        ram[176][31:0] = 32'd3483917983;
        ram[176][63:32] = 32'd27834463;
        ram[176][95:64] = 32'd2933746373;
        ram[176][127:96] = 32'd2221999411;
        ram[177][31:0] = 32'd1052551570;
        ram[177][63:32] = 32'd3550218121;
        ram[177][95:64] = 32'd140022409;
        ram[177][127:96] = 32'd1464840222;
        ram[178][31:0] = 32'd852913394;
        ram[178][63:32] = 32'd190684252;
        ram[178][95:64] = 32'd3962921086;
        ram[178][127:96] = 32'd2594523358;
        ram[179][31:0] = 32'd2485877949;
        ram[179][63:32] = 32'd486330492;
        ram[179][95:64] = 32'd47298885;
        ram[179][127:96] = 32'd3913089050;
        ram[180][31:0] = 32'd3410268326;
        ram[180][63:32] = 32'd3620424643;
        ram[180][95:64] = 32'd1996037175;
        ram[180][127:96] = 32'd485450652;
        ram[181][31:0] = 32'd705318809;
        ram[181][63:32] = 32'd3080046408;
        ram[181][95:64] = 32'd4101723380;
        ram[181][127:96] = 32'd1097647790;
        ram[182][31:0] = 32'd3542905408;
        ram[182][63:32] = 32'd1951530555;
        ram[182][95:64] = 32'd2434536837;
        ram[182][127:96] = 32'd780405641;
        ram[183][31:0] = 32'd1756047701;
        ram[183][63:32] = 32'd1592260895;
        ram[183][95:64] = 32'd1601943788;
        ram[183][127:96] = 32'd894928856;
        ram[184][31:0] = 32'd986423063;
        ram[184][63:32] = 32'd3539109186;
        ram[184][95:64] = 32'd3246599441;
        ram[184][127:96] = 32'd3879861704;
        ram[185][31:0] = 32'd1695013347;
        ram[185][63:32] = 32'd3825964589;
        ram[185][95:64] = 32'd3001673332;
        ram[185][127:96] = 32'd556542528;
        ram[186][31:0] = 32'd1702935462;
        ram[186][63:32] = 32'd824087716;
        ram[186][95:64] = 32'd1147892354;
        ram[186][127:96] = 32'd2378961500;
        ram[187][31:0] = 32'd310538191;
        ram[187][63:32] = 32'd1788156813;
        ram[187][95:64] = 32'd80903859;
        ram[187][127:96] = 32'd2915964714;
        ram[188][31:0] = 32'd2403500250;
        ram[188][63:32] = 32'd2959231921;
        ram[188][95:64] = 32'd1522336256;
        ram[188][127:96] = 32'd349850499;
        ram[189][31:0] = 32'd4214488400;
        ram[189][63:32] = 32'd3975357248;
        ram[189][95:64] = 32'd3021000205;
        ram[189][127:96] = 32'd3503267731;
        ram[190][31:0] = 32'd2429908637;
        ram[190][63:32] = 32'd3474247220;
        ram[190][95:64] = 32'd447989063;
        ram[190][127:96] = 32'd2202485930;
        ram[191][31:0] = 32'd2125336049;
        ram[191][63:32] = 32'd3634275176;
        ram[191][95:64] = 32'd2649969743;
        ram[191][127:96] = 32'd1956744276;
        ram[192][31:0] = 32'd521266459;
        ram[192][63:32] = 32'd2812677734;
        ram[192][95:64] = 32'd3061996993;
        ram[192][127:96] = 32'd1030475862;
        ram[193][31:0] = 32'd1656105210;
        ram[193][63:32] = 32'd1846218975;
        ram[193][95:64] = 32'd3672349084;
        ram[193][127:96] = 32'd515219377;
        ram[194][31:0] = 32'd2726783519;
        ram[194][63:32] = 32'd891121323;
        ram[194][95:64] = 32'd1166195020;
        ram[194][127:96] = 32'd2230018642;
        ram[195][31:0] = 32'd2527754555;
        ram[195][63:32] = 32'd1631762083;
        ram[195][95:64] = 32'd1898941484;
        ram[195][127:96] = 32'd1047929416;
        ram[196][31:0] = 32'd1886530748;
        ram[196][63:32] = 32'd1209496261;
        ram[196][95:64] = 32'd2215613352;
        ram[196][127:96] = 32'd1733548719;
        ram[197][31:0] = 32'd1647863726;
        ram[197][63:32] = 32'd1497512075;
        ram[197][95:64] = 32'd352952418;
        ram[197][127:96] = 32'd2708474774;
        ram[198][31:0] = 32'd2160729826;
        ram[198][63:32] = 32'd1811241968;
        ram[198][95:64] = 32'd3501008240;
        ram[198][127:96] = 32'd4091524596;
        ram[199][31:0] = 32'd1877609457;
        ram[199][63:32] = 32'd1827696675;
        ram[199][95:64] = 32'd3715808831;
        ram[199][127:96] = 32'd3269403007;
        ram[200][31:0] = 32'd356101764;
        ram[200][63:32] = 32'd4030133163;
        ram[200][95:64] = 32'd1172436856;
        ram[200][127:96] = 32'd3130885866;
        ram[201][31:0] = 32'd1700099309;
        ram[201][63:32] = 32'd3103250482;
        ram[201][95:64] = 32'd2394794120;
        ram[201][127:96] = 32'd3616112041;
        ram[202][31:0] = 32'd3196563487;
        ram[202][63:32] = 32'd3797926032;
        ram[202][95:64] = 32'd1249729923;
        ram[202][127:96] = 32'd3644261013;
        ram[203][31:0] = 32'd244388845;
        ram[203][63:32] = 32'd1567399322;
        ram[203][95:64] = 32'd2725263772;
        ram[203][127:96] = 32'd1145239468;
        ram[204][31:0] = 32'd3992413874;
        ram[204][63:32] = 32'd783070984;
        ram[204][95:64] = 32'd805557714;
        ram[204][127:96] = 32'd4093330237;
        ram[205][31:0] = 32'd3540865897;
        ram[205][63:32] = 32'd2641923197;
        ram[205][95:64] = 32'd2897676526;
        ram[205][127:96] = 32'd803767947;
        ram[206][31:0] = 32'd3616832036;
        ram[206][63:32] = 32'd2843325391;
        ram[206][95:64] = 32'd1511462300;
        ram[206][127:96] = 32'd3433780831;
        ram[207][31:0] = 32'd3486781950;
        ram[207][63:32] = 32'd2744509025;
        ram[207][95:64] = 32'd2106790694;
        ram[207][127:96] = 32'd2989084624;
        ram[208][31:0] = 32'd636608990;
        ram[208][63:32] = 32'd2060550887;
        ram[208][95:64] = 32'd2565041108;
        ram[208][127:96] = 32'd2346246843;
        ram[209][31:0] = 32'd374999801;
        ram[209][63:32] = 32'd2883404476;
        ram[209][95:64] = 32'd1505196816;
        ram[209][127:96] = 32'd3103203807;
        ram[210][31:0] = 32'd1961400636;
        ram[210][63:32] = 32'd1259693096;
        ram[210][95:64] = 32'd3244270472;
        ram[210][127:96] = 32'd1999149385;
        ram[211][31:0] = 32'd3760661512;
        ram[211][63:32] = 32'd2007080822;
        ram[211][95:64] = 32'd2513345585;
        ram[211][127:96] = 32'd1337120610;
        ram[212][31:0] = 32'd4157002771;
        ram[212][63:32] = 32'd1713558479;
        ram[212][95:64] = 32'd567116122;
        ram[212][127:96] = 32'd2901349547;
        ram[213][31:0] = 32'd309025837;
        ram[213][63:32] = 32'd1269596835;
        ram[213][95:64] = 32'd1000086386;
        ram[213][127:96] = 32'd3556722367;
        ram[214][31:0] = 32'd2869966604;
        ram[214][63:32] = 32'd788309353;
        ram[214][95:64] = 32'd1460621344;
        ram[214][127:96] = 32'd61833049;
        ram[215][31:0] = 32'd542097023;
        ram[215][63:32] = 32'd2384202932;
        ram[215][95:64] = 32'd2887997876;
        ram[215][127:96] = 32'd1939476593;
        ram[216][31:0] = 32'd2258396381;
        ram[216][63:32] = 32'd2384212187;
        ram[216][95:64] = 32'd2222183747;
        ram[216][127:96] = 32'd914319215;
        ram[217][31:0] = 32'd3122240770;
        ram[217][63:32] = 32'd1353029302;
        ram[217][95:64] = 32'd2534380821;
        ram[217][127:96] = 32'd2168891075;
        ram[218][31:0] = 32'd3336681769;
        ram[218][63:32] = 32'd341906945;
        ram[218][95:64] = 32'd25727163;
        ram[218][127:96] = 32'd477340108;
        ram[219][31:0] = 32'd481651494;
        ram[219][63:32] = 32'd3703124324;
        ram[219][95:64] = 32'd2455685957;
        ram[219][127:96] = 32'd1464330775;
        ram[220][31:0] = 32'd3456511089;
        ram[220][63:32] = 32'd1506016935;
        ram[220][95:64] = 32'd3835130572;
        ram[220][127:96] = 32'd3004317571;
        ram[221][31:0] = 32'd422576570;
        ram[221][63:32] = 32'd3895218455;
        ram[221][95:64] = 32'd2147679253;
        ram[221][127:96] = 32'd3092087050;
        ram[222][31:0] = 32'd309666434;
        ram[222][63:32] = 32'd955985398;
        ram[222][95:64] = 32'd3259517725;
        ram[222][127:96] = 32'd514451412;
        ram[223][31:0] = 32'd1499118016;
        ram[223][63:32] = 32'd2707802790;
        ram[223][95:64] = 32'd2339641347;
        ram[223][127:96] = 32'd653469184;
        ram[224][31:0] = 32'd1456229272;
        ram[224][63:32] = 32'd2184965099;
        ram[224][95:64] = 32'd1668711176;
        ram[224][127:96] = 32'd2631058382;
        ram[225][31:0] = 32'd2401073967;
        ram[225][63:32] = 32'd3853423062;
        ram[225][95:64] = 32'd3321083730;
        ram[225][127:96] = 32'd3146695517;
        ram[226][31:0] = 32'd365232946;
        ram[226][63:32] = 32'd1713938088;
        ram[226][95:64] = 32'd3531140847;
        ram[226][127:96] = 32'd1045330292;
        ram[227][31:0] = 32'd1536284508;
        ram[227][63:32] = 32'd1069087929;
        ram[227][95:64] = 32'd2992384195;
        ram[227][127:96] = 32'd1530098036;
        ram[228][31:0] = 32'd1888499141;
        ram[228][63:32] = 32'd714474144;
        ram[228][95:64] = 32'd3208838380;
        ram[228][127:96] = 32'd166559383;
        ram[229][31:0] = 32'd3060363333;
        ram[229][63:32] = 32'd1271364502;
        ram[229][95:64] = 32'd4239968030;
        ram[229][127:96] = 32'd1276445078;
        ram[230][31:0] = 32'd3606140741;
        ram[230][63:32] = 32'd662140256;
        ram[230][95:64] = 32'd2966286665;
        ram[230][127:96] = 32'd1827564675;
        ram[231][31:0] = 32'd605793086;
        ram[231][63:32] = 32'd164526863;
        ram[231][95:64] = 32'd2588329358;
        ram[231][127:96] = 32'd2111508981;
        ram[232][31:0] = 32'd4042835584;
        ram[232][63:32] = 32'd4115151129;
        ram[232][95:64] = 32'd3058555497;
        ram[232][127:96] = 32'd954960192;
        ram[233][31:0] = 32'd1498951355;
        ram[233][63:32] = 32'd735405892;
        ram[233][95:64] = 32'd3936725344;
        ram[233][127:96] = 32'd3119130326;
        ram[234][31:0] = 32'd1644966816;
        ram[234][63:32] = 32'd3177806684;
        ram[234][95:64] = 32'd3703155137;
        ram[234][127:96] = 32'd2577363635;
        ram[235][31:0] = 32'd3647786915;
        ram[235][63:32] = 32'd1981406870;
        ram[235][95:64] = 32'd3647750292;
        ram[235][127:96] = 32'd3360306346;
        ram[236][31:0] = 32'd1863590316;
        ram[236][63:32] = 32'd3068243404;
        ram[236][95:64] = 32'd3610640006;
        ram[236][127:96] = 32'd1282791533;
        ram[237][31:0] = 32'd3621345128;
        ram[237][63:32] = 32'd896759247;
        ram[237][95:64] = 32'd2791873980;
        ram[237][127:96] = 32'd52482036;
        ram[238][31:0] = 32'd3444183392;
        ram[238][63:32] = 32'd702849432;
        ram[238][95:64] = 32'd247955198;
        ram[238][127:96] = 32'd2403570559;
        ram[239][31:0] = 32'd3553837212;
        ram[239][63:32] = 32'd2362907167;
        ram[239][95:64] = 32'd3879054770;
        ram[239][127:96] = 32'd789581969;
        ram[240][31:0] = 32'd102932153;
        ram[240][63:32] = 32'd1879829849;
        ram[240][95:64] = 32'd3564986056;
        ram[240][127:96] = 32'd3547831979;
        ram[241][31:0] = 32'd3871364827;
        ram[241][63:32] = 32'd1400461858;
        ram[241][95:64] = 32'd3326283328;
        ram[241][127:96] = 32'd2283602290;
        ram[242][31:0] = 32'd380593856;
        ram[242][63:32] = 32'd2228588555;
        ram[242][95:64] = 32'd1184433772;
        ram[242][127:96] = 32'd2956302870;
        ram[243][31:0] = 32'd1407407298;
        ram[243][63:32] = 32'd214877909;
        ram[243][95:64] = 32'd1727455379;
        ram[243][127:96] = 32'd3749386507;
        ram[244][31:0] = 32'd3318750734;
        ram[244][63:32] = 32'd892255078;
        ram[244][95:64] = 32'd2804270651;
        ram[244][127:96] = 32'd2404684302;
        ram[245][31:0] = 32'd3450353417;
        ram[245][63:32] = 32'd377640581;
        ram[245][95:64] = 32'd3325073124;
        ram[245][127:96] = 32'd2445947169;
        ram[246][31:0] = 32'd1855044601;
        ram[246][63:32] = 32'd1066237360;
        ram[246][95:64] = 32'd1526347273;
        ram[246][127:96] = 32'd3846821607;
        ram[247][31:0] = 32'd257511150;
        ram[247][63:32] = 32'd4226538478;
        ram[247][95:64] = 32'd76974876;
        ram[247][127:96] = 32'd3252950735;
        ram[248][31:0] = 32'd3935506262;
        ram[248][63:32] = 32'd3007876411;
        ram[248][95:64] = 32'd1334459439;
        ram[248][127:96] = 32'd469208157;
        ram[249][31:0] = 32'd822061510;
        ram[249][63:32] = 32'd3817905348;
        ram[249][95:64] = 32'd876875783;
        ram[249][127:96] = 32'd3854254352;
        ram[250][31:0] = 32'd3694084155;
        ram[250][63:32] = 32'd249958146;
        ram[250][95:64] = 32'd3199440246;
        ram[250][127:96] = 32'd4260677593;
        ram[251][31:0] = 32'd1738736882;
        ram[251][63:32] = 32'd1422766232;
        ram[251][95:64] = 32'd2893698330;
        ram[251][127:96] = 32'd1819841142;
        ram[252][31:0] = 32'd2879552693;
        ram[252][63:32] = 32'd4292225377;
        ram[252][95:64] = 32'd3905914762;
        ram[252][127:96] = 32'd1770695701;
        ram[253][31:0] = 32'd3522404999;
        ram[253][63:32] = 32'd3767514378;
        ram[253][95:64] = 32'd3489533602;
        ram[253][127:96] = 32'd1511947800;
        ram[254][31:0] = 32'd1067461211;
        ram[254][63:32] = 32'd1942864530;
        ram[254][95:64] = 32'd2561367759;
        ram[254][127:96] = 32'd2891487709;
        ram[255][31:0] = 32'd1493206180;
        ram[255][63:32] = 32'd349429309;
        ram[255][95:64] = 32'd2782636993;
        ram[255][127:96] = 32'd1545197175;

    end
    always @(posedge clk) begin
        addr_r <= raddr;
        if(we) ram[waddr] <= din;
    end
    assign dout = ram[addr_r]; 

endmodule
