
/*
本文件是一个测试文件，用于测试cache模块
工作原理是模仿CPU的读写请求，对cache进行读写操作
将Cache返回的数据与预先数据进行比较，如果一致则测试通过
*/
`timescale 1ns/1ps
module cache_tb();

    //测试参数
    parameter READ_NUM = 2000;  // 测试次数 这里设置为2000次读，1000次写
    parameter WRITE_NUM = 1000;  
    //模块参数
    parameter INDEX_WIDTH       = 3;   // Cache索引位宽 2^3=8行
    parameter LINE_OFFSET_WIDTH = 2;   // 行偏移位宽，决定了一行的宽度 2^2=4字
    parameter SPACE_OFFSET      = 2;   // 一个地址空间占1个字节，因此一个字需要4个地址空间，由于假设为整字读取，处理地址的时候可以默认后两位为0
    parameter MEM_ADDR_WIDTH    = 10;   // 为了简化，这里假设内存地址宽度为10位（CPU请求地址仍然是32位，只不过我们这里简化处理，截断了高位） 
    parameter WAY_NUM           = 1;   // Cache N路组相联(N=1的时候是直接映射)

    // 变化的信号 CPU发出
    reg clk=1;
    reg rstn=1;
    reg stat=0;
    // 等rstn信号稳定后 clk信号才开始翻转
    initial begin
        #1 rstn = 0;
        #1 rstn = 1;
        stat = 1;
    end
    always  #1 clk = ~clk;

    wire [31:0] addr;
    wire r_req;
    wire w_req;
    wire [31:0] w_data;

    // 导线
    wire [31:0] r_data;
    wire miss;
    wire mem_r;
    wire mem_w;
    wire [31:0] mem_addr;
    wire [127:0] mem_w_data;
    wire [127:0] mem_r_data;
    wire mem_ready;

    // 用于测试的信号
    reg [MEM_ADDR_WIDTH-1:0] test_addr[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试地址
    reg [32:0] test_data[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试数据 最高位用于标记是否写入 0：读 1：写
    reg [31:0] test_cnt=0;  // 用于计数，每次读写操作后加1
    reg diff=0;  // 用于标记是否有不一致的数据

    // 用于对比的提交，当前cache应该给出的数据
    wire op;
    wire[31:0] data;
    assign op = test_data[test_cnt-1][32];
    assign data = test_data[test_cnt-1][31:0];
    
    // 状态机
    assign addr = test_addr[test_cnt]<<SPACE_OFFSET;
    assign r_req = test_data[test_cnt][32] == 0 ? 1 : 0;
    assign w_req = test_data[test_cnt][32] == 1 ? 1 : 0;
    assign w_data = test_data[test_cnt][31:0];
    always @(posedge clk) begin
        if (!miss && (test_cnt < READ_NUM+WRITE_NUM) && stat) begin
            if (test_data[test_cnt-1][32] == 0) begin  // 读
                if (r_data != test_data[test_cnt-1][31:0]) begin
                    $display("Read error at %d, expect %h, get %h", test_cnt, test_data[test_cnt-1][31:0], r_data);
                    diff = 1;
                end
            end
            test_cnt <= test_cnt + 1;
        end
    end

    // 例化cache
    cache #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .WAY_NUM(WAY_NUM)
    ) cache_inst(
        .clk(clk),
        .rstn(rstn),
        .addr(addr),
        .r_req(r_req),
        .w_req(w_req),
        .w_data(w_data),
        .r_data(r_data),
        .miss(miss),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 内存
    mem #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .MEM_ADDR_WIDTH(MEM_ADDR_WIDTH-LINE_OFFSET_WIDTH),
        .WAY_NUM(WAY_NUM)
    ) mem_inst(
        .clk(clk),
        .rstn(rstn),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 初始化测试数据
    initial begin
        test_addr[0] = 0;
        test_data[0] = 33'd1052567479;
        test_addr[1] = 1;
        test_data[1] = 33'd3962591981;
        test_addr[2] = 2;
        test_data[2] = 33'd5156788142;
        test_addr[3] = 905;
        test_data[3] = 33'd1713938088;
        test_addr[4] = 906;
        test_data[4] = 33'd3531140847;
        test_addr[5] = 907;
        test_data[5] = 33'd1045330292;
        test_addr[6] = 3;
        test_data[6] = 33'd7343537914;
        test_addr[7] = 4;
        test_data[7] = 33'd3294865998;
        test_addr[8] = 5;
        test_data[8] = 33'd4552824423;
        test_addr[9] = 6;
        test_data[9] = 33'd4003091934;
        test_addr[10] = 7;
        test_data[10] = 33'd3045195451;
        test_addr[11] = 8;
        test_data[11] = 33'd606447009;
        test_addr[12] = 9;
        test_data[12] = 33'd1508884471;
        test_addr[13] = 10;
        test_data[13] = 33'd4388460657;
        test_addr[14] = 11;
        test_data[14] = 33'd5997920806;
        test_addr[15] = 12;
        test_data[15] = 33'd770777372;
        test_addr[16] = 13;
        test_data[16] = 33'd675467997;
        test_addr[17] = 14;
        test_data[17] = 33'd1785532064;
        test_addr[18] = 15;
        test_data[18] = 33'd440331261;
        test_addr[19] = 16;
        test_data[19] = 33'd1426394555;
        test_addr[20] = 17;
        test_data[20] = 33'd713149634;
        test_addr[21] = 18;
        test_data[21] = 33'd3721935424;
        test_addr[22] = 19;
        test_data[22] = 33'd694124835;
        test_addr[23] = 20;
        test_data[23] = 33'd3887719615;
        test_addr[24] = 21;
        test_data[24] = 33'd6271254635;
        test_addr[25] = 22;
        test_data[25] = 33'd3582627947;
        test_addr[26] = 186;
        test_data[26] = 33'd3269096103;
        test_addr[27] = 187;
        test_data[27] = 33'd4935216646;
        test_addr[28] = 188;
        test_data[28] = 33'd3715826206;
        test_addr[29] = 189;
        test_data[29] = 33'd5424392529;
        test_addr[30] = 23;
        test_data[30] = 33'd789024827;
        test_addr[31] = 24;
        test_data[31] = 33'd6026071195;
        test_addr[32] = 25;
        test_data[32] = 33'd3096215726;
        test_addr[33] = 26;
        test_data[33] = 33'd59093393;
        test_addr[34] = 27;
        test_data[34] = 33'd1793516677;
        test_addr[35] = 28;
        test_data[35] = 33'd3711284261;
        test_addr[36] = 29;
        test_data[36] = 33'd7598114388;
        test_addr[37] = 30;
        test_data[37] = 33'd280682631;
        test_addr[38] = 31;
        test_data[38] = 33'd5647170997;
        test_addr[39] = 32;
        test_data[39] = 33'd7023115482;
        test_addr[40] = 33;
        test_data[40] = 33'd7877372138;
        test_addr[41] = 34;
        test_data[41] = 33'd3140383792;
        test_addr[42] = 35;
        test_data[42] = 33'd6118185129;
        test_addr[43] = 36;
        test_data[43] = 33'd3203529788;
        test_addr[44] = 37;
        test_data[44] = 33'd1883382384;
        test_addr[45] = 38;
        test_data[45] = 33'd5277351678;
        test_addr[46] = 39;
        test_data[46] = 33'd2778868458;
        test_addr[47] = 40;
        test_data[47] = 33'd334310572;
        test_addr[48] = 41;
        test_data[48] = 33'd5192030778;
        test_addr[49] = 42;
        test_data[49] = 33'd631245937;
        test_addr[50] = 43;
        test_data[50] = 33'd2262236211;
        test_addr[51] = 44;
        test_data[51] = 33'd2295093428;
        test_addr[52] = 45;
        test_data[52] = 33'd7760117950;
        test_addr[53] = 46;
        test_data[53] = 33'd3718565962;
        test_addr[54] = 47;
        test_data[54] = 33'd456343954;
        test_addr[55] = 211;
        test_data[55] = 33'd5525731872;
        test_addr[56] = 212;
        test_data[56] = 33'd3427452440;
        test_addr[57] = 213;
        test_data[57] = 33'd3842928591;
        test_addr[58] = 214;
        test_data[58] = 33'd67071196;
        test_addr[59] = 215;
        test_data[59] = 33'd1968456532;
        test_addr[60] = 216;
        test_data[60] = 33'd3763448983;
        test_addr[61] = 217;
        test_data[61] = 33'd91812431;
        test_addr[62] = 218;
        test_data[62] = 33'd709857341;
        test_addr[63] = 219;
        test_data[63] = 33'd6394351716;
        test_addr[64] = 220;
        test_data[64] = 33'd3956104701;
        test_addr[65] = 221;
        test_data[65] = 33'd6737584966;
        test_addr[66] = 222;
        test_data[66] = 33'd128119112;
        test_addr[67] = 223;
        test_data[67] = 33'd1645865683;
        test_addr[68] = 224;
        test_data[68] = 33'd1160411914;
        test_addr[69] = 225;
        test_data[69] = 33'd638184484;
        test_addr[70] = 226;
        test_data[70] = 33'd6428105865;
        test_addr[71] = 227;
        test_data[71] = 33'd3087655498;
        test_addr[72] = 228;
        test_data[72] = 33'd1874932830;
        test_addr[73] = 229;
        test_data[73] = 33'd5819871364;
        test_addr[74] = 230;
        test_data[74] = 33'd377097911;
        test_addr[75] = 231;
        test_data[75] = 33'd8277018722;
        test_addr[76] = 232;
        test_data[76] = 33'd4569351480;
        test_addr[77] = 233;
        test_data[77] = 33'd4982029751;
        test_addr[78] = 48;
        test_data[78] = 33'd3884411445;
        test_addr[79] = 49;
        test_data[79] = 33'd8028396518;
        test_addr[80] = 50;
        test_data[80] = 33'd4649238069;
        test_addr[81] = 51;
        test_data[81] = 33'd2846119786;
        test_addr[82] = 52;
        test_data[82] = 33'd2810219511;
        test_addr[83] = 53;
        test_data[83] = 33'd4067531662;
        test_addr[84] = 54;
        test_data[84] = 33'd1273374471;
        test_addr[85] = 55;
        test_data[85] = 33'd855085249;
        test_addr[86] = 56;
        test_data[86] = 33'd2040694399;
        test_addr[87] = 57;
        test_data[87] = 33'd3664626015;
        test_addr[88] = 58;
        test_data[88] = 33'd1265219196;
        test_addr[89] = 59;
        test_data[89] = 33'd7391994718;
        test_addr[90] = 60;
        test_data[90] = 33'd6531875140;
        test_addr[91] = 61;
        test_data[91] = 33'd468031354;
        test_addr[92] = 62;
        test_data[92] = 33'd4504848635;
        test_addr[93] = 63;
        test_data[93] = 33'd812315635;
        test_addr[94] = 64;
        test_data[94] = 33'd819283579;
        test_addr[95] = 65;
        test_data[95] = 33'd7690691796;
        test_addr[96] = 66;
        test_data[96] = 33'd2714239827;
        test_addr[97] = 67;
        test_data[97] = 33'd3494148640;
        test_addr[98] = 68;
        test_data[98] = 33'd88490023;
        test_addr[99] = 69;
        test_data[99] = 33'd2018933038;
        test_addr[100] = 70;
        test_data[100] = 33'd1396858963;
        test_addr[101] = 71;
        test_data[101] = 33'd3173125001;
        test_addr[102] = 72;
        test_data[102] = 33'd1361381559;
        test_addr[103] = 73;
        test_data[103] = 33'd546788671;
        test_addr[104] = 74;
        test_data[104] = 33'd6749477618;
        test_addr[105] = 351;
        test_data[105] = 33'd1483615543;
        test_addr[106] = 352;
        test_data[106] = 33'd6758951861;
        test_addr[107] = 353;
        test_data[107] = 33'd6792326551;
        test_addr[108] = 354;
        test_data[108] = 33'd4104199402;
        test_addr[109] = 355;
        test_data[109] = 33'd4231388117;
        test_addr[110] = 356;
        test_data[110] = 33'd328648182;
        test_addr[111] = 357;
        test_data[111] = 33'd2244387970;
        test_addr[112] = 358;
        test_data[112] = 33'd2281669903;
        test_addr[113] = 359;
        test_data[113] = 33'd4540168342;
        test_addr[114] = 360;
        test_data[114] = 33'd1685941148;
        test_addr[115] = 361;
        test_data[115] = 33'd5525071424;
        test_addr[116] = 362;
        test_data[116] = 33'd2761902832;
        test_addr[117] = 75;
        test_data[117] = 33'd1791303464;
        test_addr[118] = 76;
        test_data[118] = 33'd3925384761;
        test_addr[119] = 372;
        test_data[119] = 33'd5518166105;
        test_addr[120] = 373;
        test_data[120] = 33'd5819806658;
        test_addr[121] = 374;
        test_data[121] = 33'd276518235;
        test_addr[122] = 375;
        test_data[122] = 33'd86563587;
        test_addr[123] = 376;
        test_data[123] = 33'd2007598323;
        test_addr[124] = 377;
        test_data[124] = 33'd2225356755;
        test_addr[125] = 378;
        test_data[125] = 33'd1683535556;
        test_addr[126] = 379;
        test_data[126] = 33'd4484902977;
        test_addr[127] = 380;
        test_data[127] = 33'd2016133482;
        test_addr[128] = 381;
        test_data[128] = 33'd1644109573;
        test_addr[129] = 382;
        test_data[129] = 33'd4333113393;
        test_addr[130] = 383;
        test_data[130] = 33'd5246525281;
        test_addr[131] = 384;
        test_data[131] = 33'd1338121990;
        test_addr[132] = 385;
        test_data[132] = 33'd1312176869;
        test_addr[133] = 386;
        test_data[133] = 33'd4833973409;
        test_addr[134] = 387;
        test_data[134] = 33'd1682531476;
        test_addr[135] = 388;
        test_data[135] = 33'd4517016986;
        test_addr[136] = 389;
        test_data[136] = 33'd3581898418;
        test_addr[137] = 390;
        test_data[137] = 33'd2619734395;
        test_addr[138] = 391;
        test_data[138] = 33'd4317849461;
        test_addr[139] = 392;
        test_data[139] = 33'd4014398129;
        test_addr[140] = 393;
        test_data[140] = 33'd1253624254;
        test_addr[141] = 394;
        test_data[141] = 33'd3249060309;
        test_addr[142] = 395;
        test_data[142] = 33'd960981275;
        test_addr[143] = 396;
        test_data[143] = 33'd5998899083;
        test_addr[144] = 397;
        test_data[144] = 33'd2655648054;
        test_addr[145] = 398;
        test_data[145] = 33'd3583158237;
        test_addr[146] = 399;
        test_data[146] = 33'd1694067374;
        test_addr[147] = 400;
        test_data[147] = 33'd2624678043;
        test_addr[148] = 401;
        test_data[148] = 33'd7945980735;
        test_addr[149] = 402;
        test_data[149] = 33'd1240298673;
        test_addr[150] = 403;
        test_data[150] = 33'd1230970457;
        test_addr[151] = 404;
        test_data[151] = 33'd2974441075;
        test_addr[152] = 405;
        test_data[152] = 33'd4700635075;
        test_addr[153] = 406;
        test_data[153] = 33'd3598914984;
        test_addr[154] = 407;
        test_data[154] = 33'd6062010623;
        test_addr[155] = 408;
        test_data[155] = 33'd2708666325;
        test_addr[156] = 409;
        test_data[156] = 33'd664332654;
        test_addr[157] = 410;
        test_data[157] = 33'd2554823396;
        test_addr[158] = 411;
        test_data[158] = 33'd1912192808;
        test_addr[159] = 412;
        test_data[159] = 33'd251190816;
        test_addr[160] = 413;
        test_data[160] = 33'd42785687;
        test_addr[161] = 414;
        test_data[161] = 33'd791976254;
        test_addr[162] = 415;
        test_data[162] = 33'd3418827215;
        test_addr[163] = 416;
        test_data[163] = 33'd3371794246;
        test_addr[164] = 417;
        test_data[164] = 33'd3457950605;
        test_addr[165] = 418;
        test_data[165] = 33'd3358504200;
        test_addr[166] = 77;
        test_data[166] = 33'd3109637631;
        test_addr[167] = 983;
        test_data[167] = 33'd4548960729;
        test_addr[168] = 984;
        test_data[168] = 33'd1855044601;
        test_addr[169] = 985;
        test_data[169] = 33'd1066237360;
        test_addr[170] = 986;
        test_data[170] = 33'd1526347273;
        test_addr[171] = 987;
        test_data[171] = 33'd3846821607;
        test_addr[172] = 78;
        test_data[172] = 33'd728046435;
        test_addr[173] = 79;
        test_data[173] = 33'd5895129605;
        test_addr[174] = 80;
        test_data[174] = 33'd7500270641;
        test_addr[175] = 81;
        test_data[175] = 33'd1252273539;
        test_addr[176] = 82;
        test_data[176] = 33'd7791091190;
        test_addr[177] = 83;
        test_data[177] = 33'd4103514108;
        test_addr[178] = 84;
        test_data[178] = 33'd3678239471;
        test_addr[179] = 85;
        test_data[179] = 33'd3558159285;
        test_addr[180] = 957;
        test_data[180] = 33'd2362907167;
        test_addr[181] = 958;
        test_data[181] = 33'd3879054770;
        test_addr[182] = 959;
        test_data[182] = 33'd789581969;
        test_addr[183] = 960;
        test_data[183] = 33'd5659232848;
        test_addr[184] = 961;
        test_data[184] = 33'd1879829849;
        test_addr[185] = 962;
        test_data[185] = 33'd3564986056;
        test_addr[186] = 963;
        test_data[186] = 33'd3547831979;
        test_addr[187] = 964;
        test_data[187] = 33'd3871364827;
        test_addr[188] = 965;
        test_data[188] = 33'd1400461858;
        test_addr[189] = 86;
        test_data[189] = 33'd2026415795;
        test_addr[190] = 87;
        test_data[190] = 33'd2832515348;
        test_addr[191] = 88;
        test_data[191] = 33'd4180574515;
        test_addr[192] = 89;
        test_data[192] = 33'd777576892;
        test_addr[193] = 90;
        test_data[193] = 33'd610397100;
        test_addr[194] = 91;
        test_data[194] = 33'd1707606940;
        test_addr[195] = 92;
        test_data[195] = 33'd732174983;
        test_addr[196] = 93;
        test_data[196] = 33'd8172849913;
        test_addr[197] = 94;
        test_data[197] = 33'd4279075714;
        test_addr[198] = 95;
        test_data[198] = 33'd4186162648;
        test_addr[199] = 96;
        test_data[199] = 33'd3668307642;
        test_addr[200] = 97;
        test_data[200] = 33'd4997392963;
        test_addr[201] = 98;
        test_data[201] = 33'd2262198691;
        test_addr[202] = 99;
        test_data[202] = 33'd8030218280;
        test_addr[203] = 100;
        test_data[203] = 33'd2509988248;
        test_addr[204] = 101;
        test_data[204] = 33'd5598046868;
        test_addr[205] = 102;
        test_data[205] = 33'd7573619735;
        test_addr[206] = 103;
        test_data[206] = 33'd1753914851;
        test_addr[207] = 910;
        test_data[207] = 33'd2992384195;
        test_addr[208] = 911;
        test_data[208] = 33'd1530098036;
        test_addr[209] = 912;
        test_data[209] = 33'd1888499141;
        test_addr[210] = 913;
        test_data[210] = 33'd714474144;
        test_addr[211] = 914;
        test_data[211] = 33'd3208838380;
        test_addr[212] = 915;
        test_data[212] = 33'd166559383;
        test_addr[213] = 916;
        test_data[213] = 33'd3060363333;
        test_addr[214] = 917;
        test_data[214] = 33'd1271364502;
        test_addr[215] = 918;
        test_data[215] = 33'd4239968030;
        test_addr[216] = 919;
        test_data[216] = 33'd6334429114;
        test_addr[217] = 920;
        test_data[217] = 33'd3606140741;
        test_addr[218] = 921;
        test_data[218] = 33'd662140256;
        test_addr[219] = 104;
        test_data[219] = 33'd2137822137;
        test_addr[220] = 105;
        test_data[220] = 33'd2079086660;
        test_addr[221] = 106;
        test_data[221] = 33'd4907733251;
        test_addr[222] = 107;
        test_data[222] = 33'd2778245487;
        test_addr[223] = 108;
        test_data[223] = 33'd7227360765;
        test_addr[224] = 109;
        test_data[224] = 33'd664815512;
        test_addr[225] = 110;
        test_data[225] = 33'd3750726883;
        test_addr[226] = 757;
        test_data[226] = 33'd5706814346;
        test_addr[227] = 758;
        test_data[227] = 33'd3021000205;
        test_addr[228] = 759;
        test_data[228] = 33'd3503267731;
        test_addr[229] = 760;
        test_data[229] = 33'd2429908637;
        test_addr[230] = 761;
        test_data[230] = 33'd7737768960;
        test_addr[231] = 762;
        test_data[231] = 33'd447989063;
        test_addr[232] = 763;
        test_data[232] = 33'd2202485930;
        test_addr[233] = 764;
        test_data[233] = 33'd2125336049;
        test_addr[234] = 765;
        test_data[234] = 33'd3634275176;
        test_addr[235] = 766;
        test_data[235] = 33'd2649969743;
        test_addr[236] = 111;
        test_data[236] = 33'd2870920926;
        test_addr[237] = 112;
        test_data[237] = 33'd53516149;
        test_addr[238] = 113;
        test_data[238] = 33'd7544558860;
        test_addr[239] = 114;
        test_data[239] = 33'd574419132;
        test_addr[240] = 115;
        test_data[240] = 33'd1787837868;
        test_addr[241] = 116;
        test_data[241] = 33'd232587118;
        test_addr[242] = 117;
        test_data[242] = 33'd6679246133;
        test_addr[243] = 118;
        test_data[243] = 33'd3910724969;
        test_addr[244] = 119;
        test_data[244] = 33'd2347492591;
        test_addr[245] = 120;
        test_data[245] = 33'd3159296284;
        test_addr[246] = 121;
        test_data[246] = 33'd1116625760;
        test_addr[247] = 122;
        test_data[247] = 33'd2382385405;
        test_addr[248] = 123;
        test_data[248] = 33'd2378157637;
        test_addr[249] = 124;
        test_data[249] = 33'd6179781445;
        test_addr[250] = 125;
        test_data[250] = 33'd6380231353;
        test_addr[251] = 126;
        test_data[251] = 33'd6501560062;
        test_addr[252] = 496;
        test_data[252] = 33'd7168539293;
        test_addr[253] = 497;
        test_data[253] = 33'd253968604;
        test_addr[254] = 498;
        test_data[254] = 33'd7356876498;
        test_addr[255] = 499;
        test_data[255] = 33'd3119393922;
        test_addr[256] = 500;
        test_data[256] = 33'd5481341538;
        test_addr[257] = 501;
        test_data[257] = 33'd4273805406;
        test_addr[258] = 502;
        test_data[258] = 33'd5731145389;
        test_addr[259] = 503;
        test_data[259] = 33'd2038481495;
        test_addr[260] = 504;
        test_data[260] = 33'd1574083226;
        test_addr[261] = 505;
        test_data[261] = 33'd3731120467;
        test_addr[262] = 506;
        test_data[262] = 33'd7283148210;
        test_addr[263] = 507;
        test_data[263] = 33'd6664793892;
        test_addr[264] = 508;
        test_data[264] = 33'd3420814826;
        test_addr[265] = 509;
        test_data[265] = 33'd282828349;
        test_addr[266] = 510;
        test_data[266] = 33'd8126652940;
        test_addr[267] = 511;
        test_data[267] = 33'd667745192;
        test_addr[268] = 512;
        test_data[268] = 33'd3815785216;
        test_addr[269] = 513;
        test_data[269] = 33'd6346429545;
        test_addr[270] = 514;
        test_data[270] = 33'd7055377957;
        test_addr[271] = 515;
        test_data[271] = 33'd5053970542;
        test_addr[272] = 516;
        test_data[272] = 33'd44690167;
        test_addr[273] = 517;
        test_data[273] = 33'd8199524589;
        test_addr[274] = 127;
        test_data[274] = 33'd1861995505;
        test_addr[275] = 128;
        test_data[275] = 33'd2999443473;
        test_addr[276] = 129;
        test_data[276] = 33'd7094969221;
        test_addr[277] = 130;
        test_data[277] = 33'd1440556275;
        test_addr[278] = 131;
        test_data[278] = 33'd3900854079;
        test_addr[279] = 525;
        test_data[279] = 33'd3236712843;
        test_addr[280] = 526;
        test_data[280] = 33'd4619076371;
        test_addr[281] = 132;
        test_data[281] = 33'd1523580593;
        test_addr[282] = 133;
        test_data[282] = 33'd2214113554;
        test_addr[283] = 134;
        test_data[283] = 33'd137763915;
        test_addr[284] = 135;
        test_data[284] = 33'd5645925657;
        test_addr[285] = 572;
        test_data[285] = 33'd4628716239;
        test_addr[286] = 573;
        test_data[286] = 33'd667426504;
        test_addr[287] = 136;
        test_data[287] = 33'd796988188;
        test_addr[288] = 137;
        test_data[288] = 33'd2021339031;
        test_addr[289] = 138;
        test_data[289] = 33'd2736216411;
        test_addr[290] = 139;
        test_data[290] = 33'd932387086;
        test_addr[291] = 140;
        test_data[291] = 33'd3627393903;
        test_addr[292] = 141;
        test_data[292] = 33'd4912448088;
        test_addr[293] = 142;
        test_data[293] = 33'd662381207;
        test_addr[294] = 143;
        test_data[294] = 33'd3652162657;
        test_addr[295] = 144;
        test_data[295] = 33'd5990748232;
        test_addr[296] = 145;
        test_data[296] = 33'd3995848082;
        test_addr[297] = 146;
        test_data[297] = 33'd7219879733;
        test_addr[298] = 147;
        test_data[298] = 33'd5071552434;
        test_addr[299] = 148;
        test_data[299] = 33'd1157076026;
        test_addr[300] = 149;
        test_data[300] = 33'd3091660807;
        test_addr[301] = 150;
        test_data[301] = 33'd2857650347;
        test_addr[302] = 151;
        test_data[302] = 33'd1274566182;
        test_addr[303] = 152;
        test_data[303] = 33'd5592501431;
        test_addr[304] = 153;
        test_data[304] = 33'd3554490906;
        test_addr[305] = 154;
        test_data[305] = 33'd3756857754;
        test_addr[306] = 155;
        test_data[306] = 33'd2556299901;
        test_addr[307] = 156;
        test_data[307] = 33'd5951417504;
        test_addr[308] = 852;
        test_data[308] = 33'd309025837;
        test_addr[309] = 853;
        test_data[309] = 33'd6589782259;
        test_addr[310] = 854;
        test_data[310] = 33'd1000086386;
        test_addr[311] = 855;
        test_data[311] = 33'd3556722367;
        test_addr[312] = 856;
        test_data[312] = 33'd6537009080;
        test_addr[313] = 857;
        test_data[313] = 33'd788309353;
        test_addr[314] = 157;
        test_data[314] = 33'd295494249;
        test_addr[315] = 907;
        test_data[315] = 33'd1045330292;
        test_addr[316] = 158;
        test_data[316] = 33'd3357021415;
        test_addr[317] = 159;
        test_data[317] = 33'd885040515;
        test_addr[318] = 160;
        test_data[318] = 33'd688845184;
        test_addr[319] = 161;
        test_data[319] = 33'd1723706081;
        test_addr[320] = 162;
        test_data[320] = 33'd262508675;
        test_addr[321] = 163;
        test_data[321] = 33'd7453726228;
        test_addr[322] = 164;
        test_data[322] = 33'd10763549;
        test_addr[323] = 165;
        test_data[323] = 33'd3249592251;
        test_addr[324] = 166;
        test_data[324] = 33'd1582126961;
        test_addr[325] = 167;
        test_data[325] = 33'd3262096531;
        test_addr[326] = 939;
        test_data[326] = 33'd5184147390;
        test_addr[327] = 940;
        test_data[327] = 33'd3647786915;
        test_addr[328] = 941;
        test_data[328] = 33'd1981406870;
        test_addr[329] = 942;
        test_data[329] = 33'd6901319135;
        test_addr[330] = 943;
        test_data[330] = 33'd3360306346;
        test_addr[331] = 944;
        test_data[331] = 33'd4429138732;
        test_addr[332] = 945;
        test_data[332] = 33'd3068243404;
        test_addr[333] = 946;
        test_data[333] = 33'd6912287396;
        test_addr[334] = 947;
        test_data[334] = 33'd1282791533;
        test_addr[335] = 948;
        test_data[335] = 33'd3621345128;
        test_addr[336] = 949;
        test_data[336] = 33'd896759247;
        test_addr[337] = 168;
        test_data[337] = 33'd3104257694;
        test_addr[338] = 947;
        test_data[338] = 33'd1282791533;
        test_addr[339] = 948;
        test_data[339] = 33'd3621345128;
        test_addr[340] = 949;
        test_data[340] = 33'd8014687061;
        test_addr[341] = 950;
        test_data[341] = 33'd7297713032;
        test_addr[342] = 951;
        test_data[342] = 33'd52482036;
        test_addr[343] = 952;
        test_data[343] = 33'd3444183392;
        test_addr[344] = 953;
        test_data[344] = 33'd702849432;
        test_addr[345] = 954;
        test_data[345] = 33'd247955198;
        test_addr[346] = 955;
        test_data[346] = 33'd2403570559;
        test_addr[347] = 956;
        test_data[347] = 33'd3553837212;
        test_addr[348] = 957;
        test_data[348] = 33'd6697288910;
        test_addr[349] = 958;
        test_data[349] = 33'd3879054770;
        test_addr[350] = 959;
        test_data[350] = 33'd789581969;
        test_addr[351] = 960;
        test_data[351] = 33'd8011793532;
        test_addr[352] = 961;
        test_data[352] = 33'd7225526321;
        test_addr[353] = 962;
        test_data[353] = 33'd3564986056;
        test_addr[354] = 963;
        test_data[354] = 33'd3547831979;
        test_addr[355] = 964;
        test_data[355] = 33'd5176384803;
        test_addr[356] = 965;
        test_data[356] = 33'd1400461858;
        test_addr[357] = 169;
        test_data[357] = 33'd1157869169;
        test_addr[358] = 170;
        test_data[358] = 33'd5278097845;
        test_addr[359] = 171;
        test_data[359] = 33'd7033915995;
        test_addr[360] = 172;
        test_data[360] = 33'd909425390;
        test_addr[361] = 173;
        test_data[361] = 33'd3560746765;
        test_addr[362] = 174;
        test_data[362] = 33'd4360970199;
        test_addr[363] = 755;
        test_data[363] = 33'd5399556111;
        test_addr[364] = 756;
        test_data[364] = 33'd4214488400;
        test_addr[365] = 757;
        test_data[365] = 33'd1411847050;
        test_addr[366] = 758;
        test_data[366] = 33'd3021000205;
        test_addr[367] = 175;
        test_data[367] = 33'd5676642774;
        test_addr[368] = 176;
        test_data[368] = 33'd1240149642;
        test_addr[369] = 177;
        test_data[369] = 33'd1530014160;
        test_addr[370] = 178;
        test_data[370] = 33'd7690475394;
        test_addr[371] = 179;
        test_data[371] = 33'd2165023982;
        test_addr[372] = 180;
        test_data[372] = 33'd4349566419;
        test_addr[373] = 181;
        test_data[373] = 33'd7555096300;
        test_addr[374] = 182;
        test_data[374] = 33'd830768617;
        test_addr[375] = 183;
        test_data[375] = 33'd8043789432;
        test_addr[376] = 184;
        test_data[376] = 33'd2586566993;
        test_addr[377] = 185;
        test_data[377] = 33'd4181767754;
        test_addr[378] = 186;
        test_data[378] = 33'd3269096103;
        test_addr[379] = 187;
        test_data[379] = 33'd640249350;
        test_addr[380] = 188;
        test_data[380] = 33'd3715826206;
        test_addr[381] = 909;
        test_data[381] = 33'd1069087929;
        test_addr[382] = 910;
        test_data[382] = 33'd7971519333;
        test_addr[383] = 911;
        test_data[383] = 33'd1530098036;
        test_addr[384] = 912;
        test_data[384] = 33'd1888499141;
        test_addr[385] = 913;
        test_data[385] = 33'd714474144;
        test_addr[386] = 914;
        test_data[386] = 33'd3208838380;
        test_addr[387] = 915;
        test_data[387] = 33'd8460636591;
        test_addr[388] = 916;
        test_data[388] = 33'd3060363333;
        test_addr[389] = 917;
        test_data[389] = 33'd1271364502;
        test_addr[390] = 918;
        test_data[390] = 33'd4239968030;
        test_addr[391] = 189;
        test_data[391] = 33'd1129425233;
        test_addr[392] = 190;
        test_data[392] = 33'd1159409871;
        test_addr[393] = 191;
        test_data[393] = 33'd8038368822;
        test_addr[394] = 192;
        test_data[394] = 33'd5981779338;
        test_addr[395] = 193;
        test_data[395] = 33'd389818431;
        test_addr[396] = 194;
        test_data[396] = 33'd6195305317;
        test_addr[397] = 195;
        test_data[397] = 33'd1068866777;
        test_addr[398] = 196;
        test_data[398] = 33'd871728998;
        test_addr[399] = 197;
        test_data[399] = 33'd3233146207;
        test_addr[400] = 198;
        test_data[400] = 33'd1825329058;
        test_addr[401] = 199;
        test_data[401] = 33'd80750494;
        test_addr[402] = 200;
        test_data[402] = 33'd2827824628;
        test_addr[403] = 201;
        test_data[403] = 33'd1105729140;
        test_addr[404] = 404;
        test_data[404] = 33'd2974441075;
        test_addr[405] = 405;
        test_data[405] = 33'd7556116324;
        test_addr[406] = 406;
        test_data[406] = 33'd3598914984;
        test_addr[407] = 407;
        test_data[407] = 33'd1767043327;
        test_addr[408] = 408;
        test_data[408] = 33'd2708666325;
        test_addr[409] = 202;
        test_data[409] = 33'd1009518837;
        test_addr[410] = 203;
        test_data[410] = 33'd8362412046;
        test_addr[411] = 204;
        test_data[411] = 33'd1243827460;
        test_addr[412] = 1012;
        test_data[412] = 33'd3522404999;
        test_addr[413] = 1013;
        test_data[413] = 33'd3767514378;
        test_addr[414] = 1014;
        test_data[414] = 33'd6762745555;
        test_addr[415] = 1015;
        test_data[415] = 33'd5680405568;
        test_addr[416] = 1016;
        test_data[416] = 33'd4954872784;
        test_addr[417] = 205;
        test_data[417] = 33'd2438118847;
        test_addr[418] = 206;
        test_data[418] = 33'd4551358209;
        test_addr[419] = 207;
        test_data[419] = 33'd867306624;
        test_addr[420] = 208;
        test_data[420] = 33'd5033673891;
        test_addr[421] = 209;
        test_data[421] = 33'd8483931401;
        test_addr[422] = 210;
        test_data[422] = 33'd7276447636;
        test_addr[423] = 211;
        test_data[423] = 33'd1230764576;
        test_addr[424] = 212;
        test_data[424] = 33'd3427452440;
        test_addr[425] = 213;
        test_data[425] = 33'd3842928591;
        test_addr[426] = 214;
        test_data[426] = 33'd67071196;
        test_addr[427] = 215;
        test_data[427] = 33'd5347492977;
        test_addr[428] = 216;
        test_data[428] = 33'd3763448983;
        test_addr[429] = 217;
        test_data[429] = 33'd91812431;
        test_addr[430] = 218;
        test_data[430] = 33'd709857341;
        test_addr[431] = 328;
        test_data[431] = 33'd3264070670;
        test_addr[432] = 329;
        test_data[432] = 33'd3283575319;
        test_addr[433] = 330;
        test_data[433] = 33'd7672921207;
        test_addr[434] = 331;
        test_data[434] = 33'd4302699928;
        test_addr[435] = 332;
        test_data[435] = 33'd4698092006;
        test_addr[436] = 333;
        test_data[436] = 33'd3504452332;
        test_addr[437] = 334;
        test_data[437] = 33'd7653100462;
        test_addr[438] = 335;
        test_data[438] = 33'd459514534;
        test_addr[439] = 219;
        test_data[439] = 33'd2099384420;
        test_addr[440] = 289;
        test_data[440] = 33'd3503208650;
        test_addr[441] = 290;
        test_data[441] = 33'd193368078;
        test_addr[442] = 291;
        test_data[442] = 33'd1270361158;
        test_addr[443] = 292;
        test_data[443] = 33'd2882588279;
        test_addr[444] = 293;
        test_data[444] = 33'd7047833457;
        test_addr[445] = 294;
        test_data[445] = 33'd1462825451;
        test_addr[446] = 295;
        test_data[446] = 33'd7608401386;
        test_addr[447] = 296;
        test_data[447] = 33'd6153943196;
        test_addr[448] = 297;
        test_data[448] = 33'd1173911246;
        test_addr[449] = 298;
        test_data[449] = 33'd2569764979;
        test_addr[450] = 299;
        test_data[450] = 33'd7595161779;
        test_addr[451] = 300;
        test_data[451] = 33'd3464558724;
        test_addr[452] = 301;
        test_data[452] = 33'd4788402819;
        test_addr[453] = 302;
        test_data[453] = 33'd7624724137;
        test_addr[454] = 220;
        test_data[454] = 33'd3956104701;
        test_addr[455] = 622;
        test_data[455] = 33'd3878932875;
        test_addr[456] = 623;
        test_data[456] = 33'd1284144988;
        test_addr[457] = 624;
        test_data[457] = 33'd2824885127;
        test_addr[458] = 625;
        test_data[458] = 33'd3903890825;
        test_addr[459] = 626;
        test_data[459] = 33'd2443222463;
        test_addr[460] = 627;
        test_data[460] = 33'd207512883;
        test_addr[461] = 221;
        test_data[461] = 33'd6808137877;
        test_addr[462] = 222;
        test_data[462] = 33'd128119112;
        test_addr[463] = 223;
        test_data[463] = 33'd1645865683;
        test_addr[464] = 224;
        test_data[464] = 33'd7485774960;
        test_addr[465] = 225;
        test_data[465] = 33'd6183711781;
        test_addr[466] = 226;
        test_data[466] = 33'd2133138569;
        test_addr[467] = 227;
        test_data[467] = 33'd3087655498;
        test_addr[468] = 228;
        test_data[468] = 33'd1874932830;
        test_addr[469] = 422;
        test_data[469] = 33'd4144966284;
        test_addr[470] = 423;
        test_data[470] = 33'd4838234416;
        test_addr[471] = 424;
        test_data[471] = 33'd8554134780;
        test_addr[472] = 425;
        test_data[472] = 33'd2959861491;
        test_addr[473] = 229;
        test_data[473] = 33'd1524904068;
        test_addr[474] = 230;
        test_data[474] = 33'd377097911;
        test_addr[475] = 231;
        test_data[475] = 33'd3982051426;
        test_addr[476] = 232;
        test_data[476] = 33'd274384184;
        test_addr[477] = 233;
        test_data[477] = 33'd4607221112;
        test_addr[478] = 234;
        test_data[478] = 33'd1388060105;
        test_addr[479] = 235;
        test_data[479] = 33'd7051252711;
        test_addr[480] = 236;
        test_data[480] = 33'd2037725383;
        test_addr[481] = 237;
        test_data[481] = 33'd1838823857;
        test_addr[482] = 238;
        test_data[482] = 33'd3263906087;
        test_addr[483] = 239;
        test_data[483] = 33'd777675197;
        test_addr[484] = 240;
        test_data[484] = 33'd2405468028;
        test_addr[485] = 90;
        test_data[485] = 33'd8190272846;
        test_addr[486] = 91;
        test_data[486] = 33'd1707606940;
        test_addr[487] = 92;
        test_data[487] = 33'd8247545669;
        test_addr[488] = 93;
        test_data[488] = 33'd4388589473;
        test_addr[489] = 94;
        test_data[489] = 33'd4279075714;
        test_addr[490] = 241;
        test_data[490] = 33'd8244734788;
        test_addr[491] = 242;
        test_data[491] = 33'd4431353899;
        test_addr[492] = 243;
        test_data[492] = 33'd975543220;
        test_addr[493] = 257;
        test_data[493] = 33'd4700756776;
        test_addr[494] = 258;
        test_data[494] = 33'd2245328102;
        test_addr[495] = 259;
        test_data[495] = 33'd964259512;
        test_addr[496] = 260;
        test_data[496] = 33'd3678551605;
        test_addr[497] = 261;
        test_data[497] = 33'd1946819819;
        test_addr[498] = 262;
        test_data[498] = 33'd5713881081;
        test_addr[499] = 263;
        test_data[499] = 33'd1923525205;
        test_addr[500] = 264;
        test_data[500] = 33'd3744119204;
        test_addr[501] = 265;
        test_data[501] = 33'd4016900671;
        test_addr[502] = 266;
        test_data[502] = 33'd1955864689;
        test_addr[503] = 267;
        test_data[503] = 33'd2586515488;
        test_addr[504] = 268;
        test_data[504] = 33'd1722456956;
        test_addr[505] = 269;
        test_data[505] = 33'd8280681627;
        test_addr[506] = 270;
        test_data[506] = 33'd3591863440;
        test_addr[507] = 271;
        test_data[507] = 33'd4184036158;
        test_addr[508] = 272;
        test_data[508] = 33'd2613524396;
        test_addr[509] = 273;
        test_data[509] = 33'd4580965531;
        test_addr[510] = 274;
        test_data[510] = 33'd1993005996;
        test_addr[511] = 275;
        test_data[511] = 33'd5987230201;
        test_addr[512] = 276;
        test_data[512] = 33'd7944167454;
        test_addr[513] = 277;
        test_data[513] = 33'd2186026964;
        test_addr[514] = 278;
        test_data[514] = 33'd2738662472;
        test_addr[515] = 279;
        test_data[515] = 33'd1394720320;
        test_addr[516] = 280;
        test_data[516] = 33'd778579737;
        test_addr[517] = 281;
        test_data[517] = 33'd5881769360;
        test_addr[518] = 282;
        test_data[518] = 33'd643220710;
        test_addr[519] = 283;
        test_data[519] = 33'd6128753795;
        test_addr[520] = 284;
        test_data[520] = 33'd450921526;
        test_addr[521] = 285;
        test_data[521] = 33'd2092726877;
        test_addr[522] = 244;
        test_data[522] = 33'd1765401337;
        test_addr[523] = 245;
        test_data[523] = 33'd1169530796;
        test_addr[524] = 246;
        test_data[524] = 33'd2920595436;
        test_addr[525] = 247;
        test_data[525] = 33'd8574708850;
        test_addr[526] = 248;
        test_data[526] = 33'd7346246379;
        test_addr[527] = 249;
        test_data[527] = 33'd1695986456;
        test_addr[528] = 250;
        test_data[528] = 33'd1214633845;
        test_addr[529] = 251;
        test_data[529] = 33'd8275731799;
        test_addr[530] = 252;
        test_data[530] = 33'd6457844693;
        test_addr[531] = 805;
        test_data[531] = 33'd3103250482;
        test_addr[532] = 806;
        test_data[532] = 33'd2394794120;
        test_addr[533] = 807;
        test_data[533] = 33'd3616112041;
        test_addr[534] = 808;
        test_data[534] = 33'd3196563487;
        test_addr[535] = 809;
        test_data[535] = 33'd5390844529;
        test_addr[536] = 810;
        test_data[536] = 33'd1249729923;
        test_addr[537] = 811;
        test_data[537] = 33'd4795243738;
        test_addr[538] = 812;
        test_data[538] = 33'd6493033404;
        test_addr[539] = 813;
        test_data[539] = 33'd1567399322;
        test_addr[540] = 814;
        test_data[540] = 33'd2725263772;
        test_addr[541] = 815;
        test_data[541] = 33'd6135518878;
        test_addr[542] = 816;
        test_data[542] = 33'd6561592296;
        test_addr[543] = 817;
        test_data[543] = 33'd783070984;
        test_addr[544] = 818;
        test_data[544] = 33'd8422508264;
        test_addr[545] = 253;
        test_data[545] = 33'd3083274420;
        test_addr[546] = 254;
        test_data[546] = 33'd6438297944;
        test_addr[547] = 255;
        test_data[547] = 33'd3333567760;
        test_addr[548] = 256;
        test_data[548] = 33'd2873197191;
        test_addr[549] = 257;
        test_data[549] = 33'd405789480;
        test_addr[550] = 258;
        test_data[550] = 33'd2245328102;
        test_addr[551] = 259;
        test_data[551] = 33'd5286932626;
        test_addr[552] = 260;
        test_data[552] = 33'd7812046464;
        test_addr[553] = 261;
        test_data[553] = 33'd1946819819;
        test_addr[554] = 262;
        test_data[554] = 33'd1418913785;
        test_addr[555] = 263;
        test_data[555] = 33'd1923525205;
        test_addr[556] = 264;
        test_data[556] = 33'd3744119204;
        test_addr[557] = 265;
        test_data[557] = 33'd4016900671;
        test_addr[558] = 266;
        test_data[558] = 33'd1955864689;
        test_addr[559] = 267;
        test_data[559] = 33'd6679138310;
        test_addr[560] = 301;
        test_data[560] = 33'd493435523;
        test_addr[561] = 302;
        test_data[561] = 33'd3329756841;
        test_addr[562] = 303;
        test_data[562] = 33'd4639616666;
        test_addr[563] = 268;
        test_data[563] = 33'd1722456956;
        test_addr[564] = 269;
        test_data[564] = 33'd6165329727;
        test_addr[565] = 270;
        test_data[565] = 33'd3591863440;
        test_addr[566] = 271;
        test_data[566] = 33'd7831999982;
        test_addr[567] = 272;
        test_data[567] = 33'd4762965646;
        test_addr[568] = 273;
        test_data[568] = 33'd5967708906;
        test_addr[569] = 274;
        test_data[569] = 33'd6373642193;
        test_addr[570] = 275;
        test_data[570] = 33'd1692262905;
        test_addr[571] = 276;
        test_data[571] = 33'd3649200158;
        test_addr[572] = 277;
        test_data[572] = 33'd2186026964;
        test_addr[573] = 278;
        test_data[573] = 33'd6950975105;
        test_addr[574] = 993;
        test_data[574] = 33'd3007876411;
        test_addr[575] = 994;
        test_data[575] = 33'd4430556811;
        test_addr[576] = 995;
        test_data[576] = 33'd8128008804;
        test_addr[577] = 996;
        test_data[577] = 33'd5039003052;
        test_addr[578] = 997;
        test_data[578] = 33'd3817905348;
        test_addr[579] = 279;
        test_data[579] = 33'd7618180430;
        test_addr[580] = 280;
        test_data[580] = 33'd4812505673;
        test_addr[581] = 281;
        test_data[581] = 33'd8224744689;
        test_addr[582] = 282;
        test_data[582] = 33'd643220710;
        test_addr[583] = 283;
        test_data[583] = 33'd1833786499;
        test_addr[584] = 284;
        test_data[584] = 33'd450921526;
        test_addr[585] = 285;
        test_data[585] = 33'd7418042366;
        test_addr[586] = 286;
        test_data[586] = 33'd782042751;
        test_addr[587] = 493;
        test_data[587] = 33'd3318295190;
        test_addr[588] = 494;
        test_data[588] = 33'd2219142457;
        test_addr[589] = 495;
        test_data[589] = 33'd2985661865;
        test_addr[590] = 287;
        test_data[590] = 33'd8223176092;
        test_addr[591] = 288;
        test_data[591] = 33'd6247778810;
        test_addr[592] = 289;
        test_data[592] = 33'd3503208650;
        test_addr[593] = 290;
        test_data[593] = 33'd193368078;
        test_addr[594] = 291;
        test_data[594] = 33'd1270361158;
        test_addr[595] = 292;
        test_data[595] = 33'd6583129805;
        test_addr[596] = 293;
        test_data[596] = 33'd2752866161;
        test_addr[597] = 294;
        test_data[597] = 33'd1462825451;
        test_addr[598] = 537;
        test_data[598] = 33'd1119348756;
        test_addr[599] = 538;
        test_data[599] = 33'd5884652115;
        test_addr[600] = 539;
        test_data[600] = 33'd7481108914;
        test_addr[601] = 540;
        test_data[601] = 33'd3375317644;
        test_addr[602] = 541;
        test_data[602] = 33'd239769310;
        test_addr[603] = 542;
        test_data[603] = 33'd4367708650;
        test_addr[604] = 543;
        test_data[604] = 33'd8160207408;
        test_addr[605] = 544;
        test_data[605] = 33'd3366506315;
        test_addr[606] = 545;
        test_data[606] = 33'd2345963143;
        test_addr[607] = 546;
        test_data[607] = 33'd3228427618;
        test_addr[608] = 547;
        test_data[608] = 33'd163397476;
        test_addr[609] = 548;
        test_data[609] = 33'd1948542852;
        test_addr[610] = 549;
        test_data[610] = 33'd4281859846;
        test_addr[611] = 550;
        test_data[611] = 33'd3804497467;
        test_addr[612] = 551;
        test_data[612] = 33'd5900690673;
        test_addr[613] = 552;
        test_data[613] = 33'd822192939;
        test_addr[614] = 553;
        test_data[614] = 33'd4863041004;
        test_addr[615] = 554;
        test_data[615] = 33'd279679526;
        test_addr[616] = 555;
        test_data[616] = 33'd3894035056;
        test_addr[617] = 556;
        test_data[617] = 33'd4546315113;
        test_addr[618] = 557;
        test_data[618] = 33'd3787715714;
        test_addr[619] = 558;
        test_data[619] = 33'd4516560427;
        test_addr[620] = 559;
        test_data[620] = 33'd3250198723;
        test_addr[621] = 560;
        test_data[621] = 33'd3966735267;
        test_addr[622] = 561;
        test_data[622] = 33'd4675864130;
        test_addr[623] = 562;
        test_data[623] = 33'd4874861904;
        test_addr[624] = 563;
        test_data[624] = 33'd2283251439;
        test_addr[625] = 564;
        test_data[625] = 33'd7800636892;
        test_addr[626] = 565;
        test_data[626] = 33'd1424860412;
        test_addr[627] = 566;
        test_data[627] = 33'd4203930147;
        test_addr[628] = 567;
        test_data[628] = 33'd6291993177;
        test_addr[629] = 568;
        test_data[629] = 33'd74969035;
        test_addr[630] = 569;
        test_data[630] = 33'd3416048394;
        test_addr[631] = 570;
        test_data[631] = 33'd3977968930;
        test_addr[632] = 571;
        test_data[632] = 33'd7835124221;
        test_addr[633] = 572;
        test_data[633] = 33'd333748943;
        test_addr[634] = 573;
        test_data[634] = 33'd667426504;
        test_addr[635] = 574;
        test_data[635] = 33'd277213762;
        test_addr[636] = 575;
        test_data[636] = 33'd2498279954;
        test_addr[637] = 576;
        test_data[637] = 33'd8295214957;
        test_addr[638] = 577;
        test_data[638] = 33'd474077448;
        test_addr[639] = 578;
        test_data[639] = 33'd2578797357;
        test_addr[640] = 579;
        test_data[640] = 33'd2429845848;
        test_addr[641] = 295;
        test_data[641] = 33'd3313434090;
        test_addr[642] = 296;
        test_data[642] = 33'd1858975900;
        test_addr[643] = 371;
        test_data[643] = 33'd4633103161;
        test_addr[644] = 372;
        test_data[644] = 33'd7137866315;
        test_addr[645] = 373;
        test_data[645] = 33'd1524839362;
        test_addr[646] = 374;
        test_data[646] = 33'd7891999687;
        test_addr[647] = 375;
        test_data[647] = 33'd86563587;
        test_addr[648] = 376;
        test_data[648] = 33'd2007598323;
        test_addr[649] = 377;
        test_data[649] = 33'd2225356755;
        test_addr[650] = 378;
        test_data[650] = 33'd1683535556;
        test_addr[651] = 379;
        test_data[651] = 33'd189935681;
        test_addr[652] = 297;
        test_data[652] = 33'd5550535678;
        test_addr[653] = 298;
        test_data[653] = 33'd5649789836;
        test_addr[654] = 567;
        test_data[654] = 33'd1997025881;
        test_addr[655] = 299;
        test_data[655] = 33'd6268728660;
        test_addr[656] = 300;
        test_data[656] = 33'd3464558724;
        test_addr[657] = 301;
        test_data[657] = 33'd493435523;
        test_addr[658] = 302;
        test_data[658] = 33'd3329756841;
        test_addr[659] = 303;
        test_data[659] = 33'd6690420131;
        test_addr[660] = 304;
        test_data[660] = 33'd3131755163;
        test_addr[661] = 305;
        test_data[661] = 33'd2985268612;
        test_addr[662] = 306;
        test_data[662] = 33'd2048220064;
        test_addr[663] = 307;
        test_data[663] = 33'd395268976;
        test_addr[664] = 308;
        test_data[664] = 33'd1555365123;
        test_addr[665] = 309;
        test_data[665] = 33'd1157989693;
        test_addr[666] = 310;
        test_data[666] = 33'd892285550;
        test_addr[667] = 311;
        test_data[667] = 33'd757719279;
        test_addr[668] = 312;
        test_data[668] = 33'd5876477841;
        test_addr[669] = 313;
        test_data[669] = 33'd2709848361;
        test_addr[670] = 314;
        test_data[670] = 33'd4792863700;
        test_addr[671] = 315;
        test_data[671] = 33'd5833393492;
        test_addr[672] = 316;
        test_data[672] = 33'd2469986364;
        test_addr[673] = 317;
        test_data[673] = 33'd1975671844;
        test_addr[674] = 318;
        test_data[674] = 33'd3064576727;
        test_addr[675] = 319;
        test_data[675] = 33'd3883511213;
        test_addr[676] = 500;
        test_data[676] = 33'd1186374242;
        test_addr[677] = 501;
        test_data[677] = 33'd7403902751;
        test_addr[678] = 320;
        test_data[678] = 33'd2659365932;
        test_addr[679] = 321;
        test_data[679] = 33'd2227829365;
        test_addr[680] = 322;
        test_data[680] = 33'd6828888674;
        test_addr[681] = 323;
        test_data[681] = 33'd200882046;
        test_addr[682] = 324;
        test_data[682] = 33'd2565321190;
        test_addr[683] = 325;
        test_data[683] = 33'd2573803079;
        test_addr[684] = 326;
        test_data[684] = 33'd4237884957;
        test_addr[685] = 327;
        test_data[685] = 33'd7226486472;
        test_addr[686] = 328;
        test_data[686] = 33'd3264070670;
        test_addr[687] = 329;
        test_data[687] = 33'd3283575319;
        test_addr[688] = 330;
        test_data[688] = 33'd3377953911;
        test_addr[689] = 331;
        test_data[689] = 33'd7732632;
        test_addr[690] = 332;
        test_data[690] = 33'd403124710;
        test_addr[691] = 333;
        test_data[691] = 33'd3504452332;
        test_addr[692] = 334;
        test_data[692] = 33'd7136595493;
        test_addr[693] = 335;
        test_data[693] = 33'd4836406072;
        test_addr[694] = 336;
        test_data[694] = 33'd966779298;
        test_addr[695] = 745;
        test_data[695] = 33'd824087716;
        test_addr[696] = 746;
        test_data[696] = 33'd1147892354;
        test_addr[697] = 747;
        test_data[697] = 33'd5034975190;
        test_addr[698] = 337;
        test_data[698] = 33'd4218420959;
        test_addr[699] = 338;
        test_data[699] = 33'd2832891657;
        test_addr[700] = 380;
        test_data[700] = 33'd5226745734;
        test_addr[701] = 381;
        test_data[701] = 33'd6025088853;
        test_addr[702] = 382;
        test_data[702] = 33'd5724345560;
        test_addr[703] = 383;
        test_data[703] = 33'd951557985;
        test_addr[704] = 339;
        test_data[704] = 33'd3901609669;
        test_addr[705] = 340;
        test_data[705] = 33'd2309224711;
        test_addr[706] = 341;
        test_data[706] = 33'd1297508340;
        test_addr[707] = 342;
        test_data[707] = 33'd3867550255;
        test_addr[708] = 343;
        test_data[708] = 33'd6937468559;
        test_addr[709] = 344;
        test_data[709] = 33'd100362266;
        test_addr[710] = 662;
        test_data[710] = 33'd6772296886;
        test_addr[711] = 663;
        test_data[711] = 33'd372966818;
        test_addr[712] = 664;
        test_data[712] = 33'd6132108558;
        test_addr[713] = 665;
        test_data[713] = 33'd4823700786;
        test_addr[714] = 666;
        test_data[714] = 33'd4072192775;
        test_addr[715] = 667;
        test_data[715] = 33'd2563820725;
        test_addr[716] = 668;
        test_data[716] = 33'd3382879701;
        test_addr[717] = 669;
        test_data[717] = 33'd3165934849;
        test_addr[718] = 670;
        test_data[718] = 33'd2503869172;
        test_addr[719] = 671;
        test_data[719] = 33'd222714301;
        test_addr[720] = 345;
        test_data[720] = 33'd2316252777;
        test_addr[721] = 346;
        test_data[721] = 33'd2418381156;
        test_addr[722] = 347;
        test_data[722] = 33'd3975745931;
        test_addr[723] = 348;
        test_data[723] = 33'd2859983252;
        test_addr[724] = 349;
        test_data[724] = 33'd2089693596;
        test_addr[725] = 350;
        test_data[725] = 33'd1993790010;
        test_addr[726] = 351;
        test_data[726] = 33'd1483615543;
        test_addr[727] = 352;
        test_data[727] = 33'd7680306837;
        test_addr[728] = 353;
        test_data[728] = 33'd2497359255;
        test_addr[729] = 354;
        test_data[729] = 33'd4104199402;
        test_addr[730] = 355;
        test_data[730] = 33'd5398725571;
        test_addr[731] = 356;
        test_data[731] = 33'd328648182;
        test_addr[732] = 357;
        test_data[732] = 33'd8276786891;
        test_addr[733] = 358;
        test_data[733] = 33'd2281669903;
        test_addr[734] = 359;
        test_data[734] = 33'd245201046;
        test_addr[735] = 360;
        test_data[735] = 33'd1685941148;
        test_addr[736] = 361;
        test_data[736] = 33'd1230104128;
        test_addr[737] = 362;
        test_data[737] = 33'd2761902832;
        test_addr[738] = 363;
        test_data[738] = 33'd803716268;
        test_addr[739] = 364;
        test_data[739] = 33'd3270560608;
        test_addr[740] = 365;
        test_data[740] = 33'd92649394;
        test_addr[741] = 366;
        test_data[741] = 33'd4105913331;
        test_addr[742] = 367;
        test_data[742] = 33'd3378755930;
        test_addr[743] = 368;
        test_data[743] = 33'd7502139528;
        test_addr[744] = 369;
        test_data[744] = 33'd2921962052;
        test_addr[745] = 552;
        test_data[745] = 33'd5774456499;
        test_addr[746] = 553;
        test_data[746] = 33'd568073708;
        test_addr[747] = 370;
        test_data[747] = 33'd1101997953;
        test_addr[748] = 371;
        test_data[748] = 33'd338135865;
        test_addr[749] = 372;
        test_data[749] = 33'd8201970068;
        test_addr[750] = 373;
        test_data[750] = 33'd1524839362;
        test_addr[751] = 374;
        test_data[751] = 33'd3597032391;
        test_addr[752] = 375;
        test_data[752] = 33'd86563587;
        test_addr[753] = 376;
        test_data[753] = 33'd2007598323;
        test_addr[754] = 377;
        test_data[754] = 33'd6864750829;
        test_addr[755] = 378;
        test_data[755] = 33'd1683535556;
        test_addr[756] = 379;
        test_data[756] = 33'd5985026329;
        test_addr[757] = 380;
        test_data[757] = 33'd931778438;
        test_addr[758] = 381;
        test_data[758] = 33'd1730121557;
        test_addr[759] = 382;
        test_data[759] = 33'd7630803241;
        test_addr[760] = 383;
        test_data[760] = 33'd4346540679;
        test_addr[761] = 384;
        test_data[761] = 33'd1338121990;
        test_addr[762] = 385;
        test_data[762] = 33'd7044698085;
        test_addr[763] = 644;
        test_data[763] = 33'd3042117089;
        test_addr[764] = 645;
        test_data[764] = 33'd3539970854;
        test_addr[765] = 646;
        test_data[765] = 33'd8296645476;
        test_addr[766] = 647;
        test_data[766] = 33'd3098822722;
        test_addr[767] = 648;
        test_data[767] = 33'd320726234;
        test_addr[768] = 649;
        test_data[768] = 33'd2831991724;
        test_addr[769] = 650;
        test_data[769] = 33'd3593391115;
        test_addr[770] = 651;
        test_data[770] = 33'd6723127522;
        test_addr[771] = 652;
        test_data[771] = 33'd5186879897;
        test_addr[772] = 653;
        test_data[772] = 33'd2986341452;
        test_addr[773] = 654;
        test_data[773] = 33'd266085065;
        test_addr[774] = 655;
        test_data[774] = 33'd763025037;
        test_addr[775] = 656;
        test_data[775] = 33'd5051010472;
        test_addr[776] = 657;
        test_data[776] = 33'd668982047;
        test_addr[777] = 658;
        test_data[777] = 33'd2565372091;
        test_addr[778] = 659;
        test_data[778] = 33'd1343443381;
        test_addr[779] = 660;
        test_data[779] = 33'd8464711346;
        test_addr[780] = 661;
        test_data[780] = 33'd5323330305;
        test_addr[781] = 662;
        test_data[781] = 33'd7409917304;
        test_addr[782] = 663;
        test_data[782] = 33'd8304218084;
        test_addr[783] = 664;
        test_data[783] = 33'd1837141262;
        test_addr[784] = 665;
        test_data[784] = 33'd6792175769;
        test_addr[785] = 666;
        test_data[785] = 33'd6192224370;
        test_addr[786] = 386;
        test_data[786] = 33'd539006113;
        test_addr[787] = 387;
        test_data[787] = 33'd1682531476;
        test_addr[788] = 388;
        test_data[788] = 33'd222049690;
        test_addr[789] = 389;
        test_data[789] = 33'd8575367807;
        test_addr[790] = 390;
        test_data[790] = 33'd2619734395;
        test_addr[791] = 391;
        test_data[791] = 33'd22882165;
        test_addr[792] = 518;
        test_data[792] = 33'd4343951664;
        test_addr[793] = 519;
        test_data[793] = 33'd1574109177;
        test_addr[794] = 392;
        test_data[794] = 33'd6749306979;
        test_addr[795] = 393;
        test_data[795] = 33'd7531889498;
        test_addr[796] = 394;
        test_data[796] = 33'd3249060309;
        test_addr[797] = 395;
        test_data[797] = 33'd4396110102;
        test_addr[798] = 928;
        test_data[798] = 33'd4042835584;
        test_addr[799] = 929;
        test_data[799] = 33'd4115151129;
        test_addr[800] = 930;
        test_data[800] = 33'd3058555497;
        test_addr[801] = 931;
        test_data[801] = 33'd4302895425;
        test_addr[802] = 932;
        test_data[802] = 33'd1498951355;
        test_addr[803] = 933;
        test_data[803] = 33'd4536004200;
        test_addr[804] = 934;
        test_data[804] = 33'd3936725344;
        test_addr[805] = 935;
        test_data[805] = 33'd3119130326;
        test_addr[806] = 936;
        test_data[806] = 33'd4988848755;
        test_addr[807] = 937;
        test_data[807] = 33'd3177806684;
        test_addr[808] = 938;
        test_data[808] = 33'd3703155137;
        test_addr[809] = 939;
        test_data[809] = 33'd889180094;
        test_addr[810] = 940;
        test_data[810] = 33'd4507518110;
        test_addr[811] = 941;
        test_data[811] = 33'd1981406870;
        test_addr[812] = 942;
        test_data[812] = 33'd2606351839;
        test_addr[813] = 396;
        test_data[813] = 33'd8002451475;
        test_addr[814] = 397;
        test_data[814] = 33'd7275093251;
        test_addr[815] = 398;
        test_data[815] = 33'd3583158237;
        test_addr[816] = 399;
        test_data[816] = 33'd1694067374;
        test_addr[817] = 400;
        test_data[817] = 33'd2624678043;
        test_addr[818] = 401;
        test_data[818] = 33'd3651013439;
        test_addr[819] = 402;
        test_data[819] = 33'd1240298673;
        test_addr[820] = 53;
        test_data[820] = 33'd5394474912;
        test_addr[821] = 54;
        test_data[821] = 33'd6907486484;
        test_addr[822] = 55;
        test_data[822] = 33'd855085249;
        test_addr[823] = 56;
        test_data[823] = 33'd2040694399;
        test_addr[824] = 57;
        test_data[824] = 33'd7473814280;
        test_addr[825] = 58;
        test_data[825] = 33'd1265219196;
        test_addr[826] = 59;
        test_data[826] = 33'd3097027422;
        test_addr[827] = 60;
        test_data[827] = 33'd4417070254;
        test_addr[828] = 61;
        test_data[828] = 33'd468031354;
        test_addr[829] = 62;
        test_data[829] = 33'd209881339;
        test_addr[830] = 403;
        test_data[830] = 33'd5115395963;
        test_addr[831] = 404;
        test_data[831] = 33'd2974441075;
        test_addr[832] = 405;
        test_data[832] = 33'd3261149028;
        test_addr[833] = 724;
        test_data[833] = 33'd7360840813;
        test_addr[834] = 725;
        test_data[834] = 33'd8526315959;
        test_addr[835] = 726;
        test_data[835] = 33'd4101723380;
        test_addr[836] = 406;
        test_data[836] = 33'd3598914984;
        test_addr[837] = 407;
        test_data[837] = 33'd1767043327;
        test_addr[838] = 408;
        test_data[838] = 33'd2708666325;
        test_addr[839] = 259;
        test_data[839] = 33'd8083756326;
        test_addr[840] = 260;
        test_data[840] = 33'd3517079168;
        test_addr[841] = 261;
        test_data[841] = 33'd1946819819;
        test_addr[842] = 262;
        test_data[842] = 33'd8115131983;
        test_addr[843] = 409;
        test_data[843] = 33'd664332654;
        test_addr[844] = 410;
        test_data[844] = 33'd2554823396;
        test_addr[845] = 411;
        test_data[845] = 33'd1912192808;
        test_addr[846] = 1004;
        test_data[846] = 33'd1738736882;
        test_addr[847] = 1005;
        test_data[847] = 33'd1422766232;
        test_addr[848] = 1006;
        test_data[848] = 33'd2893698330;
        test_addr[849] = 1007;
        test_data[849] = 33'd1819841142;
        test_addr[850] = 1008;
        test_data[850] = 33'd2879552693;
        test_addr[851] = 1009;
        test_data[851] = 33'd4292225377;
        test_addr[852] = 1010;
        test_data[852] = 33'd3905914762;
        test_addr[853] = 1011;
        test_data[853] = 33'd1770695701;
        test_addr[854] = 1012;
        test_data[854] = 33'd3522404999;
        test_addr[855] = 1013;
        test_data[855] = 33'd7062350654;
        test_addr[856] = 1014;
        test_data[856] = 33'd2467778259;
        test_addr[857] = 1015;
        test_data[857] = 33'd1385438272;
        test_addr[858] = 1016;
        test_data[858] = 33'd659905488;
        test_addr[859] = 412;
        test_data[859] = 33'd5431733346;
        test_addr[860] = 413;
        test_data[860] = 33'd42785687;
        test_addr[861] = 414;
        test_data[861] = 33'd4945397945;
        test_addr[862] = 415;
        test_data[862] = 33'd3418827215;
        test_addr[863] = 416;
        test_data[863] = 33'd3371794246;
        test_addr[864] = 629;
        test_data[864] = 33'd3640747;
        test_addr[865] = 630;
        test_data[865] = 33'd2440170518;
        test_addr[866] = 631;
        test_data[866] = 33'd243801277;
        test_addr[867] = 632;
        test_data[867] = 33'd6979379595;
        test_addr[868] = 633;
        test_data[868] = 33'd3766781495;
        test_addr[869] = 634;
        test_data[869] = 33'd941110408;
        test_addr[870] = 417;
        test_data[870] = 33'd7904599271;
        test_addr[871] = 418;
        test_data[871] = 33'd4735005430;
        test_addr[872] = 419;
        test_data[872] = 33'd3137721503;
        test_addr[873] = 420;
        test_data[873] = 33'd3236855211;
        test_addr[874] = 421;
        test_data[874] = 33'd5044363472;
        test_addr[875] = 422;
        test_data[875] = 33'd4144966284;
        test_addr[876] = 423;
        test_data[876] = 33'd543267120;
        test_addr[877] = 424;
        test_data[877] = 33'd4259167484;
        test_addr[878] = 425;
        test_data[878] = 33'd2959861491;
        test_addr[879] = 426;
        test_data[879] = 33'd4113724443;
        test_addr[880] = 427;
        test_data[880] = 33'd3990194643;
        test_addr[881] = 457;
        test_data[881] = 33'd2500934454;
        test_addr[882] = 458;
        test_data[882] = 33'd2264632454;
        test_addr[883] = 459;
        test_data[883] = 33'd8099435533;
        test_addr[884] = 460;
        test_data[884] = 33'd2220856156;
        test_addr[885] = 461;
        test_data[885] = 33'd3428994727;
        test_addr[886] = 462;
        test_data[886] = 33'd4446020023;
        test_addr[887] = 463;
        test_data[887] = 33'd6015469463;
        test_addr[888] = 464;
        test_data[888] = 33'd8390278337;
        test_addr[889] = 465;
        test_data[889] = 33'd3508624685;
        test_addr[890] = 466;
        test_data[890] = 33'd6055986827;
        test_addr[891] = 467;
        test_data[891] = 33'd1066574642;
        test_addr[892] = 468;
        test_data[892] = 33'd1244655582;
        test_addr[893] = 469;
        test_data[893] = 33'd4275884649;
        test_addr[894] = 470;
        test_data[894] = 33'd1434334882;
        test_addr[895] = 471;
        test_data[895] = 33'd3824336063;
        test_addr[896] = 472;
        test_data[896] = 33'd4261511285;
        test_addr[897] = 473;
        test_data[897] = 33'd3858581669;
        test_addr[898] = 474;
        test_data[898] = 33'd4537685587;
        test_addr[899] = 428;
        test_data[899] = 33'd3112127436;
        test_addr[900] = 96;
        test_data[900] = 33'd7340107857;
        test_addr[901] = 97;
        test_data[901] = 33'd702425667;
        test_addr[902] = 98;
        test_data[902] = 33'd2262198691;
        test_addr[903] = 99;
        test_data[903] = 33'd3735250984;
        test_addr[904] = 100;
        test_data[904] = 33'd2509988248;
        test_addr[905] = 101;
        test_data[905] = 33'd1303079572;
        test_addr[906] = 102;
        test_data[906] = 33'd7027788573;
        test_addr[907] = 429;
        test_data[907] = 33'd4791663874;
        test_addr[908] = 430;
        test_data[908] = 33'd3912201120;
        test_addr[909] = 431;
        test_data[909] = 33'd6379223070;
        test_addr[910] = 432;
        test_data[910] = 33'd807161466;
        test_addr[911] = 433;
        test_data[911] = 33'd363795349;
        test_addr[912] = 434;
        test_data[912] = 33'd7293721338;
        test_addr[913] = 435;
        test_data[913] = 33'd2035856504;
        test_addr[914] = 436;
        test_data[914] = 33'd8568290205;
        test_addr[915] = 437;
        test_data[915] = 33'd1332405155;
        test_addr[916] = 438;
        test_data[916] = 33'd6460754832;
        test_addr[917] = 439;
        test_data[917] = 33'd1956260871;
        test_addr[918] = 440;
        test_data[918] = 33'd2562872072;
        test_addr[919] = 552;
        test_data[919] = 33'd5355052870;
        test_addr[920] = 553;
        test_data[920] = 33'd568073708;
        test_addr[921] = 554;
        test_data[921] = 33'd5259500731;
        test_addr[922] = 555;
        test_data[922] = 33'd3894035056;
        test_addr[923] = 556;
        test_data[923] = 33'd251347817;
        test_addr[924] = 557;
        test_data[924] = 33'd7656331289;
        test_addr[925] = 558;
        test_data[925] = 33'd221593131;
        test_addr[926] = 559;
        test_data[926] = 33'd3250198723;
        test_addr[927] = 560;
        test_data[927] = 33'd3966735267;
        test_addr[928] = 561;
        test_data[928] = 33'd5372436028;
        test_addr[929] = 562;
        test_data[929] = 33'd579894608;
        test_addr[930] = 563;
        test_data[930] = 33'd2283251439;
        test_addr[931] = 564;
        test_data[931] = 33'd3505669596;
        test_addr[932] = 565;
        test_data[932] = 33'd5271239953;
        test_addr[933] = 566;
        test_data[933] = 33'd4203930147;
        test_addr[934] = 567;
        test_data[934] = 33'd1997025881;
        test_addr[935] = 568;
        test_data[935] = 33'd74969035;
        test_addr[936] = 569;
        test_data[936] = 33'd3416048394;
        test_addr[937] = 570;
        test_data[937] = 33'd3977968930;
        test_addr[938] = 441;
        test_data[938] = 33'd65904936;
        test_addr[939] = 442;
        test_data[939] = 33'd1741314760;
        test_addr[940] = 443;
        test_data[940] = 33'd5371030409;
        test_addr[941] = 444;
        test_data[941] = 33'd4084632541;
        test_addr[942] = 445;
        test_data[942] = 33'd3196251038;
        test_addr[943] = 446;
        test_data[943] = 33'd6763356948;
        test_addr[944] = 447;
        test_data[944] = 33'd7610765084;
        test_addr[945] = 448;
        test_data[945] = 33'd1265298441;
        test_addr[946] = 449;
        test_data[946] = 33'd2908833870;
        test_addr[947] = 450;
        test_data[947] = 33'd2162667854;
        test_addr[948] = 872;
        test_data[948] = 33'd5620553560;
        test_addr[949] = 873;
        test_data[949] = 33'd6691719662;
        test_addr[950] = 874;
        test_data[950] = 33'd25727163;
        test_addr[951] = 875;
        test_data[951] = 33'd477340108;
        test_addr[952] = 876;
        test_data[952] = 33'd5606990723;
        test_addr[953] = 877;
        test_data[953] = 33'd3703124324;
        test_addr[954] = 878;
        test_data[954] = 33'd7378662421;
        test_addr[955] = 879;
        test_data[955] = 33'd1464330775;
        test_addr[956] = 880;
        test_data[956] = 33'd4549146278;
        test_addr[957] = 451;
        test_data[957] = 33'd7782778936;
        test_addr[958] = 452;
        test_data[958] = 33'd8011060688;
        test_addr[959] = 453;
        test_data[959] = 33'd285543293;
        test_addr[960] = 454;
        test_data[960] = 33'd2191347482;
        test_addr[961] = 455;
        test_data[961] = 33'd2580577157;
        test_addr[962] = 456;
        test_data[962] = 33'd321448812;
        test_addr[963] = 457;
        test_data[963] = 33'd2500934454;
        test_addr[964] = 458;
        test_data[964] = 33'd2264632454;
        test_addr[965] = 459;
        test_data[965] = 33'd3804468237;
        test_addr[966] = 460;
        test_data[966] = 33'd2220856156;
        test_addr[967] = 461;
        test_data[967] = 33'd3428994727;
        test_addr[968] = 462;
        test_data[968] = 33'd151052727;
        test_addr[969] = 463;
        test_data[969] = 33'd1720502167;
        test_addr[970] = 464;
        test_data[970] = 33'd6120160395;
        test_addr[971] = 465;
        test_data[971] = 33'd3508624685;
        test_addr[972] = 466;
        test_data[972] = 33'd1761019531;
        test_addr[973] = 467;
        test_data[973] = 33'd1066574642;
        test_addr[974] = 468;
        test_data[974] = 33'd4843926671;
        test_addr[975] = 469;
        test_data[975] = 33'd4275884649;
        test_addr[976] = 470;
        test_data[976] = 33'd1434334882;
        test_addr[977] = 419;
        test_data[977] = 33'd3137721503;
        test_addr[978] = 420;
        test_data[978] = 33'd4412783747;
        test_addr[979] = 471;
        test_data[979] = 33'd3824336063;
        test_addr[980] = 899;
        test_data[980] = 33'd2631058382;
        test_addr[981] = 472;
        test_data[981] = 33'd4468450433;
        test_addr[982] = 473;
        test_data[982] = 33'd3858581669;
        test_addr[983] = 474;
        test_data[983] = 33'd242718291;
        test_addr[984] = 475;
        test_data[984] = 33'd3328634438;
        test_addr[985] = 476;
        test_data[985] = 33'd2866816344;
        test_addr[986] = 477;
        test_data[986] = 33'd3782855187;
        test_addr[987] = 478;
        test_data[987] = 33'd6437917831;
        test_addr[988] = 755;
        test_data[988] = 33'd1104588815;
        test_addr[989] = 756;
        test_data[989] = 33'd7842182917;
        test_addr[990] = 479;
        test_data[990] = 33'd6588385089;
        test_addr[991] = 480;
        test_data[991] = 33'd799026300;
        test_addr[992] = 481;
        test_data[992] = 33'd3611509395;
        test_addr[993] = 364;
        test_data[993] = 33'd3270560608;
        test_addr[994] = 365;
        test_data[994] = 33'd4719062742;
        test_addr[995] = 366;
        test_data[995] = 33'd4105913331;
        test_addr[996] = 367;
        test_data[996] = 33'd3378755930;
        test_addr[997] = 368;
        test_data[997] = 33'd3207172232;
        test_addr[998] = 369;
        test_data[998] = 33'd2921962052;
        test_addr[999] = 370;
        test_data[999] = 33'd1101997953;
        test_addr[1000] = 371;
        test_data[1000] = 33'd338135865;
        test_addr[1001] = 372;
        test_data[1001] = 33'd4900288633;
        test_addr[1002] = 373;
        test_data[1002] = 33'd1524839362;
        test_addr[1003] = 482;
        test_data[1003] = 33'd4402868585;
        test_addr[1004] = 754;
        test_data[1004] = 33'd1522336256;
        test_addr[1005] = 755;
        test_data[1005] = 33'd1104588815;
        test_addr[1006] = 756;
        test_data[1006] = 33'd5342596311;
        test_addr[1007] = 757;
        test_data[1007] = 33'd1411847050;
        test_addr[1008] = 483;
        test_data[1008] = 33'd3314459181;
        test_addr[1009] = 484;
        test_data[1009] = 33'd5093760048;
        test_addr[1010] = 485;
        test_data[1010] = 33'd453359906;
        test_addr[1011] = 486;
        test_data[1011] = 33'd8188830353;
        test_addr[1012] = 487;
        test_data[1012] = 33'd7953507360;
        test_addr[1013] = 488;
        test_data[1013] = 33'd1111823230;
        test_addr[1014] = 489;
        test_data[1014] = 33'd1327010194;
        test_addr[1015] = 490;
        test_data[1015] = 33'd1847146603;
        test_addr[1016] = 491;
        test_data[1016] = 33'd6649522250;
        test_addr[1017] = 492;
        test_data[1017] = 33'd2825740953;
        test_addr[1018] = 493;
        test_data[1018] = 33'd8418113341;
        test_addr[1019] = 494;
        test_data[1019] = 33'd2219142457;
        test_addr[1020] = 495;
        test_data[1020] = 33'd6902331883;
        test_addr[1021] = 496;
        test_data[1021] = 33'd7263515245;
        test_addr[1022] = 497;
        test_data[1022] = 33'd253968604;
        test_addr[1023] = 498;
        test_data[1023] = 33'd3061909202;
        test_addr[1024] = 499;
        test_data[1024] = 33'd6106764415;
        test_addr[1025] = 500;
        test_data[1025] = 33'd1186374242;
        test_addr[1026] = 501;
        test_data[1026] = 33'd7019881564;
        test_addr[1027] = 1017;
        test_data[1027] = 33'd1942864530;
        test_addr[1028] = 1018;
        test_data[1028] = 33'd6014433002;
        test_addr[1029] = 1019;
        test_data[1029] = 33'd2891487709;
        test_addr[1030] = 1020;
        test_data[1030] = 33'd1493206180;
        test_addr[1031] = 502;
        test_data[1031] = 33'd6377533717;
        test_addr[1032] = 503;
        test_data[1032] = 33'd7229823078;
        test_addr[1033] = 504;
        test_data[1033] = 33'd1574083226;
        test_addr[1034] = 189;
        test_data[1034] = 33'd5261376945;
        test_addr[1035] = 190;
        test_data[1035] = 33'd1159409871;
        test_addr[1036] = 191;
        test_data[1036] = 33'd3743401526;
        test_addr[1037] = 192;
        test_data[1037] = 33'd1686812042;
        test_addr[1038] = 193;
        test_data[1038] = 33'd389818431;
        test_addr[1039] = 194;
        test_data[1039] = 33'd5882511768;
        test_addr[1040] = 195;
        test_data[1040] = 33'd1068866777;
        test_addr[1041] = 505;
        test_data[1041] = 33'd3731120467;
        test_addr[1042] = 506;
        test_data[1042] = 33'd2988180914;
        test_addr[1043] = 507;
        test_data[1043] = 33'd6060339491;
        test_addr[1044] = 508;
        test_data[1044] = 33'd3420814826;
        test_addr[1045] = 509;
        test_data[1045] = 33'd282828349;
        test_addr[1046] = 510;
        test_data[1046] = 33'd3831685644;
        test_addr[1047] = 511;
        test_data[1047] = 33'd667745192;
        test_addr[1048] = 919;
        test_data[1048] = 33'd2039461818;
        test_addr[1049] = 920;
        test_data[1049] = 33'd3606140741;
        test_addr[1050] = 921;
        test_data[1050] = 33'd662140256;
        test_addr[1051] = 922;
        test_data[1051] = 33'd2966286665;
        test_addr[1052] = 923;
        test_data[1052] = 33'd1827564675;
        test_addr[1053] = 924;
        test_data[1053] = 33'd605793086;
        test_addr[1054] = 512;
        test_data[1054] = 33'd6106755207;
        test_addr[1055] = 513;
        test_data[1055] = 33'd2051462249;
        test_addr[1056] = 514;
        test_data[1056] = 33'd2760410661;
        test_addr[1057] = 515;
        test_data[1057] = 33'd7637287168;
        test_addr[1058] = 516;
        test_data[1058] = 33'd7179112593;
        test_addr[1059] = 517;
        test_data[1059] = 33'd4457231055;
        test_addr[1060] = 518;
        test_data[1060] = 33'd48984368;
        test_addr[1061] = 519;
        test_data[1061] = 33'd1574109177;
        test_addr[1062] = 520;
        test_data[1062] = 33'd847712690;
        test_addr[1063] = 521;
        test_data[1063] = 33'd8381387186;
        test_addr[1064] = 522;
        test_data[1064] = 33'd4674569930;
        test_addr[1065] = 523;
        test_data[1065] = 33'd40985424;
        test_addr[1066] = 524;
        test_data[1066] = 33'd3607396520;
        test_addr[1067] = 525;
        test_data[1067] = 33'd3236712843;
        test_addr[1068] = 526;
        test_data[1068] = 33'd324109075;
        test_addr[1069] = 527;
        test_data[1069] = 33'd7495486352;
        test_addr[1070] = 528;
        test_data[1070] = 33'd5617230810;
        test_addr[1071] = 529;
        test_data[1071] = 33'd1798434561;
        test_addr[1072] = 530;
        test_data[1072] = 33'd7866367211;
        test_addr[1073] = 531;
        test_data[1073] = 33'd1917508662;
        test_addr[1074] = 532;
        test_data[1074] = 33'd7570608729;
        test_addr[1075] = 180;
        test_data[1075] = 33'd54599123;
        test_addr[1076] = 181;
        test_data[1076] = 33'd3260129004;
        test_addr[1077] = 182;
        test_data[1077] = 33'd830768617;
        test_addr[1078] = 183;
        test_data[1078] = 33'd5113234577;
        test_addr[1079] = 184;
        test_data[1079] = 33'd2586566993;
        test_addr[1080] = 185;
        test_data[1080] = 33'd4181767754;
        test_addr[1081] = 186;
        test_data[1081] = 33'd3269096103;
        test_addr[1082] = 187;
        test_data[1082] = 33'd640249350;
        test_addr[1083] = 188;
        test_data[1083] = 33'd7596521115;
        test_addr[1084] = 189;
        test_data[1084] = 33'd966409649;
        test_addr[1085] = 533;
        test_data[1085] = 33'd5264424910;
        test_addr[1086] = 275;
        test_data[1086] = 33'd1692262905;
        test_addr[1087] = 276;
        test_data[1087] = 33'd5926162428;
        test_addr[1088] = 277;
        test_data[1088] = 33'd2186026964;
        test_addr[1089] = 278;
        test_data[1089] = 33'd5271386823;
        test_addr[1090] = 279;
        test_data[1090] = 33'd3323213134;
        test_addr[1091] = 280;
        test_data[1091] = 33'd517538377;
        test_addr[1092] = 281;
        test_data[1092] = 33'd3929777393;
        test_addr[1093] = 282;
        test_data[1093] = 33'd643220710;
        test_addr[1094] = 283;
        test_data[1094] = 33'd1833786499;
        test_addr[1095] = 284;
        test_data[1095] = 33'd5603055021;
        test_addr[1096] = 285;
        test_data[1096] = 33'd4849316648;
        test_addr[1097] = 286;
        test_data[1097] = 33'd6489874367;
        test_addr[1098] = 287;
        test_data[1098] = 33'd3928208796;
        test_addr[1099] = 288;
        test_data[1099] = 33'd1952811514;
        test_addr[1100] = 289;
        test_data[1100] = 33'd3503208650;
        test_addr[1101] = 290;
        test_data[1101] = 33'd193368078;
        test_addr[1102] = 291;
        test_data[1102] = 33'd1270361158;
        test_addr[1103] = 292;
        test_data[1103] = 33'd2288162509;
        test_addr[1104] = 293;
        test_data[1104] = 33'd6098839160;
        test_addr[1105] = 294;
        test_data[1105] = 33'd1462825451;
        test_addr[1106] = 534;
        test_data[1106] = 33'd7609099576;
        test_addr[1107] = 535;
        test_data[1107] = 33'd740792702;
        test_addr[1108] = 536;
        test_data[1108] = 33'd1359838887;
        test_addr[1109] = 537;
        test_data[1109] = 33'd1119348756;
        test_addr[1110] = 538;
        test_data[1110] = 33'd8274520020;
        test_addr[1111] = 539;
        test_data[1111] = 33'd3186141618;
        test_addr[1112] = 540;
        test_data[1112] = 33'd4587297326;
        test_addr[1113] = 541;
        test_data[1113] = 33'd239769310;
        test_addr[1114] = 542;
        test_data[1114] = 33'd72741354;
        test_addr[1115] = 543;
        test_data[1115] = 33'd7684069834;
        test_addr[1116] = 544;
        test_data[1116] = 33'd3366506315;
        test_addr[1117] = 545;
        test_data[1117] = 33'd2345963143;
        test_addr[1118] = 546;
        test_data[1118] = 33'd3228427618;
        test_addr[1119] = 547;
        test_data[1119] = 33'd8446464250;
        test_addr[1120] = 548;
        test_data[1120] = 33'd5467155352;
        test_addr[1121] = 549;
        test_data[1121] = 33'd8018311090;
        test_addr[1122] = 550;
        test_data[1122] = 33'd3804497467;
        test_addr[1123] = 551;
        test_data[1123] = 33'd8104880645;
        test_addr[1124] = 552;
        test_data[1124] = 33'd8056299463;
        test_addr[1125] = 553;
        test_data[1125] = 33'd568073708;
        test_addr[1126] = 554;
        test_data[1126] = 33'd964533435;
        test_addr[1127] = 555;
        test_data[1127] = 33'd3894035056;
        test_addr[1128] = 86;
        test_data[1128] = 33'd7673239827;
        test_addr[1129] = 87;
        test_data[1129] = 33'd2832515348;
        test_addr[1130] = 88;
        test_data[1130] = 33'd5756290695;
        test_addr[1131] = 89;
        test_data[1131] = 33'd777576892;
        test_addr[1132] = 90;
        test_data[1132] = 33'd3895305550;
        test_addr[1133] = 556;
        test_data[1133] = 33'd251347817;
        test_addr[1134] = 557;
        test_data[1134] = 33'd5612825308;
        test_addr[1135] = 558;
        test_data[1135] = 33'd221593131;
        test_addr[1136] = 559;
        test_data[1136] = 33'd8553918342;
        test_addr[1137] = 560;
        test_data[1137] = 33'd8302946213;
        test_addr[1138] = 561;
        test_data[1138] = 33'd1077468732;
        test_addr[1139] = 562;
        test_data[1139] = 33'd579894608;
        test_addr[1140] = 563;
        test_data[1140] = 33'd2283251439;
        test_addr[1141] = 564;
        test_data[1141] = 33'd7229791127;
        test_addr[1142] = 565;
        test_data[1142] = 33'd976272657;
        test_addr[1143] = 566;
        test_data[1143] = 33'd7611456480;
        test_addr[1144] = 567;
        test_data[1144] = 33'd1997025881;
        test_addr[1145] = 568;
        test_data[1145] = 33'd74969035;
        test_addr[1146] = 902;
        test_data[1146] = 33'd3321083730;
        test_addr[1147] = 903;
        test_data[1147] = 33'd3146695517;
        test_addr[1148] = 904;
        test_data[1148] = 33'd7067277155;
        test_addr[1149] = 905;
        test_data[1149] = 33'd1713938088;
        test_addr[1150] = 906;
        test_data[1150] = 33'd3531140847;
        test_addr[1151] = 907;
        test_data[1151] = 33'd1045330292;
        test_addr[1152] = 908;
        test_data[1152] = 33'd6471499310;
        test_addr[1153] = 909;
        test_data[1153] = 33'd1069087929;
        test_addr[1154] = 910;
        test_data[1154] = 33'd3676552037;
        test_addr[1155] = 911;
        test_data[1155] = 33'd4579493945;
        test_addr[1156] = 912;
        test_data[1156] = 33'd1888499141;
        test_addr[1157] = 913;
        test_data[1157] = 33'd714474144;
        test_addr[1158] = 914;
        test_data[1158] = 33'd6270762888;
        test_addr[1159] = 915;
        test_data[1159] = 33'd4165669295;
        test_addr[1160] = 916;
        test_data[1160] = 33'd3060363333;
        test_addr[1161] = 917;
        test_data[1161] = 33'd5478774957;
        test_addr[1162] = 918;
        test_data[1162] = 33'd4239968030;
        test_addr[1163] = 919;
        test_data[1163] = 33'd7025860956;
        test_addr[1164] = 569;
        test_data[1164] = 33'd5047719948;
        test_addr[1165] = 570;
        test_data[1165] = 33'd3977968930;
        test_addr[1166] = 497;
        test_data[1166] = 33'd4300685245;
        test_addr[1167] = 498;
        test_data[1167] = 33'd8588315097;
        test_addr[1168] = 499;
        test_data[1168] = 33'd6101537607;
        test_addr[1169] = 500;
        test_data[1169] = 33'd1186374242;
        test_addr[1170] = 501;
        test_data[1170] = 33'd2724914268;
        test_addr[1171] = 502;
        test_data[1171] = 33'd6917074800;
        test_addr[1172] = 503;
        test_data[1172] = 33'd4833786369;
        test_addr[1173] = 571;
        test_data[1173] = 33'd3540156925;
        test_addr[1174] = 572;
        test_data[1174] = 33'd8171889624;
        test_addr[1175] = 573;
        test_data[1175] = 33'd667426504;
        test_addr[1176] = 574;
        test_data[1176] = 33'd277213762;
        test_addr[1177] = 575;
        test_data[1177] = 33'd7340152710;
        test_addr[1178] = 576;
        test_data[1178] = 33'd4000247661;
        test_addr[1179] = 577;
        test_data[1179] = 33'd474077448;
        test_addr[1180] = 578;
        test_data[1180] = 33'd2578797357;
        test_addr[1181] = 330;
        test_data[1181] = 33'd3377953911;
        test_addr[1182] = 331;
        test_data[1182] = 33'd7732632;
        test_addr[1183] = 332;
        test_data[1183] = 33'd403124710;
        test_addr[1184] = 333;
        test_data[1184] = 33'd3504452332;
        test_addr[1185] = 334;
        test_data[1185] = 33'd2841628197;
        test_addr[1186] = 335;
        test_data[1186] = 33'd6521233655;
        test_addr[1187] = 336;
        test_data[1187] = 33'd5040289745;
        test_addr[1188] = 337;
        test_data[1188] = 33'd4218420959;
        test_addr[1189] = 338;
        test_data[1189] = 33'd2832891657;
        test_addr[1190] = 339;
        test_data[1190] = 33'd7532254382;
        test_addr[1191] = 340;
        test_data[1191] = 33'd2309224711;
        test_addr[1192] = 341;
        test_data[1192] = 33'd1297508340;
        test_addr[1193] = 342;
        test_data[1193] = 33'd3867550255;
        test_addr[1194] = 343;
        test_data[1194] = 33'd2642501263;
        test_addr[1195] = 344;
        test_data[1195] = 33'd100362266;
        test_addr[1196] = 345;
        test_data[1196] = 33'd4379718114;
        test_addr[1197] = 346;
        test_data[1197] = 33'd2418381156;
        test_addr[1198] = 347;
        test_data[1198] = 33'd6682985408;
        test_addr[1199] = 348;
        test_data[1199] = 33'd2859983252;
        test_addr[1200] = 579;
        test_data[1200] = 33'd6518911936;
        test_addr[1201] = 580;
        test_data[1201] = 33'd3083515047;
        test_addr[1202] = 581;
        test_data[1202] = 33'd7204371839;
        test_addr[1203] = 262;
        test_data[1203] = 33'd7905717909;
        test_addr[1204] = 263;
        test_data[1204] = 33'd5292915570;
        test_addr[1205] = 264;
        test_data[1205] = 33'd4542373727;
        test_addr[1206] = 265;
        test_data[1206] = 33'd4016900671;
        test_addr[1207] = 266;
        test_data[1207] = 33'd1955864689;
        test_addr[1208] = 267;
        test_data[1208] = 33'd2384171014;
        test_addr[1209] = 268;
        test_data[1209] = 33'd8430857312;
        test_addr[1210] = 269;
        test_data[1210] = 33'd1870362431;
        test_addr[1211] = 270;
        test_data[1211] = 33'd3591863440;
        test_addr[1212] = 271;
        test_data[1212] = 33'd5676684663;
        test_addr[1213] = 272;
        test_data[1213] = 33'd5827929463;
        test_addr[1214] = 273;
        test_data[1214] = 33'd1672741610;
        test_addr[1215] = 274;
        test_data[1215] = 33'd2078674897;
        test_addr[1216] = 275;
        test_data[1216] = 33'd7021143707;
        test_addr[1217] = 276;
        test_data[1217] = 33'd6883287131;
        test_addr[1218] = 582;
        test_data[1218] = 33'd2220997705;
        test_addr[1219] = 200;
        test_data[1219] = 33'd2827824628;
        test_addr[1220] = 201;
        test_data[1220] = 33'd7675494397;
        test_addr[1221] = 202;
        test_data[1221] = 33'd5542347112;
        test_addr[1222] = 203;
        test_data[1222] = 33'd7919769411;
        test_addr[1223] = 583;
        test_data[1223] = 33'd2367557065;
        test_addr[1224] = 584;
        test_data[1224] = 33'd4897203055;
        test_addr[1225] = 504;
        test_data[1225] = 33'd1574083226;
        test_addr[1226] = 505;
        test_data[1226] = 33'd3731120467;
        test_addr[1227] = 506;
        test_data[1227] = 33'd2988180914;
        test_addr[1228] = 507;
        test_data[1228] = 33'd1765372195;
        test_addr[1229] = 585;
        test_data[1229] = 33'd3545634013;
        test_addr[1230] = 586;
        test_data[1230] = 33'd3351735354;
        test_addr[1231] = 587;
        test_data[1231] = 33'd291280601;
        test_addr[1232] = 588;
        test_data[1232] = 33'd6318957505;
        test_addr[1233] = 589;
        test_data[1233] = 33'd5618684185;
        test_addr[1234] = 590;
        test_data[1234] = 33'd4931530400;
        test_addr[1235] = 745;
        test_data[1235] = 33'd5728956167;
        test_addr[1236] = 746;
        test_data[1236] = 33'd7303851618;
        test_addr[1237] = 747;
        test_data[1237] = 33'd740007894;
        test_addr[1238] = 748;
        test_data[1238] = 33'd310538191;
        test_addr[1239] = 591;
        test_data[1239] = 33'd4103338995;
        test_addr[1240] = 592;
        test_data[1240] = 33'd3890705901;
        test_addr[1241] = 593;
        test_data[1241] = 33'd58166058;
        test_addr[1242] = 594;
        test_data[1242] = 33'd8420808485;
        test_addr[1243] = 595;
        test_data[1243] = 33'd8031590255;
        test_addr[1244] = 596;
        test_data[1244] = 33'd3005148523;
        test_addr[1245] = 597;
        test_data[1245] = 33'd3336186297;
        test_addr[1246] = 598;
        test_data[1246] = 33'd4433093745;
        test_addr[1247] = 79;
        test_data[1247] = 33'd7858842824;
        test_addr[1248] = 80;
        test_data[1248] = 33'd3205303345;
        test_addr[1249] = 81;
        test_data[1249] = 33'd1252273539;
        test_addr[1250] = 82;
        test_data[1250] = 33'd3496123894;
        test_addr[1251] = 83;
        test_data[1251] = 33'd5360081232;
        test_addr[1252] = 84;
        test_data[1252] = 33'd3678239471;
        test_addr[1253] = 85;
        test_data[1253] = 33'd3558159285;
        test_addr[1254] = 86;
        test_data[1254] = 33'd3378272531;
        test_addr[1255] = 87;
        test_data[1255] = 33'd7258027848;
        test_addr[1256] = 88;
        test_data[1256] = 33'd1461323399;
        test_addr[1257] = 89;
        test_data[1257] = 33'd777576892;
        test_addr[1258] = 90;
        test_data[1258] = 33'd3895305550;
        test_addr[1259] = 91;
        test_data[1259] = 33'd1707606940;
        test_addr[1260] = 92;
        test_data[1260] = 33'd4537437257;
        test_addr[1261] = 93;
        test_data[1261] = 33'd93622177;
        test_addr[1262] = 94;
        test_data[1262] = 33'd4279075714;
        test_addr[1263] = 95;
        test_data[1263] = 33'd4186162648;
        test_addr[1264] = 96;
        test_data[1264] = 33'd5809815071;
        test_addr[1265] = 97;
        test_data[1265] = 33'd702425667;
        test_addr[1266] = 98;
        test_data[1266] = 33'd6482254222;
        test_addr[1267] = 99;
        test_data[1267] = 33'd8196413094;
        test_addr[1268] = 100;
        test_data[1268] = 33'd5509561754;
        test_addr[1269] = 101;
        test_data[1269] = 33'd1303079572;
        test_addr[1270] = 102;
        test_data[1270] = 33'd2732821277;
        test_addr[1271] = 103;
        test_data[1271] = 33'd1753914851;
        test_addr[1272] = 104;
        test_data[1272] = 33'd2137822137;
        test_addr[1273] = 599;
        test_data[1273] = 33'd7905633535;
        test_addr[1274] = 600;
        test_data[1274] = 33'd508264472;
        test_addr[1275] = 601;
        test_data[1275] = 33'd2571072663;
        test_addr[1276] = 602;
        test_data[1276] = 33'd2987575655;
        test_addr[1277] = 678;
        test_data[1277] = 33'd2364391312;
        test_addr[1278] = 679;
        test_data[1278] = 33'd5713521064;
        test_addr[1279] = 680;
        test_data[1279] = 33'd708134854;
        test_addr[1280] = 681;
        test_data[1280] = 33'd2488012861;
        test_addr[1281] = 682;
        test_data[1281] = 33'd2655148014;
        test_addr[1282] = 683;
        test_data[1282] = 33'd3868012904;
        test_addr[1283] = 603;
        test_data[1283] = 33'd6675343823;
        test_addr[1284] = 604;
        test_data[1284] = 33'd1222723850;
        test_addr[1285] = 605;
        test_data[1285] = 33'd3919297631;
        test_addr[1286] = 606;
        test_data[1286] = 33'd242612497;
        test_addr[1287] = 607;
        test_data[1287] = 33'd7304109004;
        test_addr[1288] = 618;
        test_data[1288] = 33'd7083904914;
        test_addr[1289] = 608;
        test_data[1289] = 33'd4136444716;
        test_addr[1290] = 609;
        test_data[1290] = 33'd3925486970;
        test_addr[1291] = 610;
        test_data[1291] = 33'd3603903628;
        test_addr[1292] = 399;
        test_data[1292] = 33'd1694067374;
        test_addr[1293] = 400;
        test_data[1293] = 33'd2624678043;
        test_addr[1294] = 401;
        test_data[1294] = 33'd3651013439;
        test_addr[1295] = 402;
        test_data[1295] = 33'd1240298673;
        test_addr[1296] = 403;
        test_data[1296] = 33'd820428667;
        test_addr[1297] = 404;
        test_data[1297] = 33'd2974441075;
        test_addr[1298] = 405;
        test_data[1298] = 33'd3261149028;
        test_addr[1299] = 406;
        test_data[1299] = 33'd3598914984;
        test_addr[1300] = 407;
        test_data[1300] = 33'd6254539809;
        test_addr[1301] = 408;
        test_data[1301] = 33'd2708666325;
        test_addr[1302] = 409;
        test_data[1302] = 33'd664332654;
        test_addr[1303] = 410;
        test_data[1303] = 33'd2554823396;
        test_addr[1304] = 411;
        test_data[1304] = 33'd1912192808;
        test_addr[1305] = 412;
        test_data[1305] = 33'd1136766050;
        test_addr[1306] = 413;
        test_data[1306] = 33'd42785687;
        test_addr[1307] = 414;
        test_data[1307] = 33'd650430649;
        test_addr[1308] = 415;
        test_data[1308] = 33'd3418827215;
        test_addr[1309] = 416;
        test_data[1309] = 33'd4324041238;
        test_addr[1310] = 417;
        test_data[1310] = 33'd3609631975;
        test_addr[1311] = 418;
        test_data[1311] = 33'd440038134;
        test_addr[1312] = 419;
        test_data[1312] = 33'd3137721503;
        test_addr[1313] = 420;
        test_data[1313] = 33'd5410495330;
        test_addr[1314] = 421;
        test_data[1314] = 33'd749396176;
        test_addr[1315] = 422;
        test_data[1315] = 33'd8424371424;
        test_addr[1316] = 423;
        test_data[1316] = 33'd543267120;
        test_addr[1317] = 611;
        test_data[1317] = 33'd2389840076;
        test_addr[1318] = 612;
        test_data[1318] = 33'd1075777044;
        test_addr[1319] = 613;
        test_data[1319] = 33'd2147567015;
        test_addr[1320] = 614;
        test_data[1320] = 33'd2943240457;
        test_addr[1321] = 615;
        test_data[1321] = 33'd2283134385;
        test_addr[1322] = 616;
        test_data[1322] = 33'd5640958638;
        test_addr[1323] = 617;
        test_data[1323] = 33'd5274421218;
        test_addr[1324] = 618;
        test_data[1324] = 33'd2788937618;
        test_addr[1325] = 619;
        test_data[1325] = 33'd3667454584;
        test_addr[1326] = 620;
        test_data[1326] = 33'd2816982930;
        test_addr[1327] = 621;
        test_data[1327] = 33'd3470453698;
        test_addr[1328] = 341;
        test_data[1328] = 33'd1297508340;
        test_addr[1329] = 622;
        test_data[1329] = 33'd3878932875;
        test_addr[1330] = 623;
        test_data[1330] = 33'd1284144988;
        test_addr[1331] = 624;
        test_data[1331] = 33'd2824885127;
        test_addr[1332] = 625;
        test_data[1332] = 33'd7538014277;
        test_addr[1333] = 701;
        test_data[1333] = 33'd2591022462;
        test_addr[1334] = 626;
        test_data[1334] = 33'd2443222463;
        test_addr[1335] = 627;
        test_data[1335] = 33'd6636608881;
        test_addr[1336] = 628;
        test_data[1336] = 33'd390612325;
        test_addr[1337] = 629;
        test_data[1337] = 33'd3640747;
        test_addr[1338] = 630;
        test_data[1338] = 33'd2440170518;
        test_addr[1339] = 631;
        test_data[1339] = 33'd243801277;
        test_addr[1340] = 632;
        test_data[1340] = 33'd6859443872;
        test_addr[1341] = 633;
        test_data[1341] = 33'd5211041330;
        test_addr[1342] = 634;
        test_data[1342] = 33'd7329083725;
        test_addr[1343] = 635;
        test_data[1343] = 33'd2142044604;
        test_addr[1344] = 342;
        test_data[1344] = 33'd3867550255;
        test_addr[1345] = 343;
        test_data[1345] = 33'd2642501263;
        test_addr[1346] = 344;
        test_data[1346] = 33'd100362266;
        test_addr[1347] = 636;
        test_data[1347] = 33'd3358336986;
        test_addr[1348] = 637;
        test_data[1348] = 33'd7746659701;
        test_addr[1349] = 638;
        test_data[1349] = 33'd2786119313;
        test_addr[1350] = 2;
        test_data[1350] = 33'd7036036440;
        test_addr[1351] = 3;
        test_data[1351] = 33'd3048570618;
        test_addr[1352] = 4;
        test_data[1352] = 33'd6848074264;
        test_addr[1353] = 5;
        test_data[1353] = 33'd5433778074;
        test_addr[1354] = 6;
        test_data[1354] = 33'd4003091934;
        test_addr[1355] = 7;
        test_data[1355] = 33'd3045195451;
        test_addr[1356] = 8;
        test_data[1356] = 33'd606447009;
        test_addr[1357] = 9;
        test_data[1357] = 33'd1508884471;
        test_addr[1358] = 10;
        test_data[1358] = 33'd93493361;
        test_addr[1359] = 11;
        test_data[1359] = 33'd5360836092;
        test_addr[1360] = 12;
        test_data[1360] = 33'd770777372;
        test_addr[1361] = 13;
        test_data[1361] = 33'd675467997;
        test_addr[1362] = 14;
        test_data[1362] = 33'd1785532064;
        test_addr[1363] = 15;
        test_data[1363] = 33'd5756267892;
        test_addr[1364] = 639;
        test_data[1364] = 33'd7935463702;
        test_addr[1365] = 640;
        test_data[1365] = 33'd1294707516;
        test_addr[1366] = 641;
        test_data[1366] = 33'd263459559;
        test_addr[1367] = 970;
        test_data[1367] = 33'd1184433772;
        test_addr[1368] = 971;
        test_data[1368] = 33'd2956302870;
        test_addr[1369] = 972;
        test_data[1369] = 33'd1407407298;
        test_addr[1370] = 973;
        test_data[1370] = 33'd214877909;
        test_addr[1371] = 974;
        test_data[1371] = 33'd1727455379;
        test_addr[1372] = 975;
        test_data[1372] = 33'd3749386507;
        test_addr[1373] = 976;
        test_data[1373] = 33'd3318750734;
        test_addr[1374] = 977;
        test_data[1374] = 33'd892255078;
        test_addr[1375] = 978;
        test_data[1375] = 33'd2804270651;
        test_addr[1376] = 979;
        test_data[1376] = 33'd4779712395;
        test_addr[1377] = 980;
        test_data[1377] = 33'd8427158991;
        test_addr[1378] = 981;
        test_data[1378] = 33'd7931822166;
        test_addr[1379] = 982;
        test_data[1379] = 33'd3325073124;
        test_addr[1380] = 983;
        test_data[1380] = 33'd253993433;
        test_addr[1381] = 984;
        test_data[1381] = 33'd1855044601;
        test_addr[1382] = 985;
        test_data[1382] = 33'd1066237360;
        test_addr[1383] = 642;
        test_data[1383] = 33'd6955893670;
        test_addr[1384] = 447;
        test_data[1384] = 33'd3315797788;
        test_addr[1385] = 448;
        test_data[1385] = 33'd1265298441;
        test_addr[1386] = 449;
        test_data[1386] = 33'd2908833870;
        test_addr[1387] = 450;
        test_data[1387] = 33'd2162667854;
        test_addr[1388] = 451;
        test_data[1388] = 33'd3487811640;
        test_addr[1389] = 452;
        test_data[1389] = 33'd4843807922;
        test_addr[1390] = 453;
        test_data[1390] = 33'd285543293;
        test_addr[1391] = 454;
        test_data[1391] = 33'd5590560255;
        test_addr[1392] = 643;
        test_data[1392] = 33'd2925530671;
        test_addr[1393] = 644;
        test_data[1393] = 33'd8253592696;
        test_addr[1394] = 645;
        test_data[1394] = 33'd3539970854;
        test_addr[1395] = 646;
        test_data[1395] = 33'd4001678180;
        test_addr[1396] = 647;
        test_data[1396] = 33'd7652880563;
        test_addr[1397] = 648;
        test_data[1397] = 33'd320726234;
        test_addr[1398] = 649;
        test_data[1398] = 33'd2831991724;
        test_addr[1399] = 650;
        test_data[1399] = 33'd3593391115;
        test_addr[1400] = 651;
        test_data[1400] = 33'd2428160226;
        test_addr[1401] = 652;
        test_data[1401] = 33'd891912601;
        test_addr[1402] = 653;
        test_data[1402] = 33'd2986341452;
        test_addr[1403] = 654;
        test_data[1403] = 33'd8274407193;
        test_addr[1404] = 655;
        test_data[1404] = 33'd763025037;
        test_addr[1405] = 656;
        test_data[1405] = 33'd756043176;
        test_addr[1406] = 657;
        test_data[1406] = 33'd668982047;
        test_addr[1407] = 658;
        test_data[1407] = 33'd2565372091;
        test_addr[1408] = 659;
        test_data[1408] = 33'd7644348422;
        test_addr[1409] = 698;
        test_data[1409] = 33'd4345694941;
        test_addr[1410] = 699;
        test_data[1410] = 33'd507075352;
        test_addr[1411] = 700;
        test_data[1411] = 33'd1049995550;
        test_addr[1412] = 701;
        test_data[1412] = 33'd2591022462;
        test_addr[1413] = 702;
        test_data[1413] = 33'd2452957524;
        test_addr[1414] = 703;
        test_data[1414] = 33'd2083865596;
        test_addr[1415] = 704;
        test_data[1415] = 33'd3483917983;
        test_addr[1416] = 705;
        test_data[1416] = 33'd27834463;
        test_addr[1417] = 706;
        test_data[1417] = 33'd6011559468;
        test_addr[1418] = 660;
        test_data[1418] = 33'd4169744050;
        test_addr[1419] = 661;
        test_data[1419] = 33'd4703301226;
        test_addr[1420] = 662;
        test_data[1420] = 33'd7877626317;
        test_addr[1421] = 663;
        test_data[1421] = 33'd5768702542;
        test_addr[1422] = 664;
        test_data[1422] = 33'd5484878242;
        test_addr[1423] = 979;
        test_data[1423] = 33'd7671727475;
        test_addr[1424] = 980;
        test_data[1424] = 33'd4132191695;
        test_addr[1425] = 981;
        test_data[1425] = 33'd3636854870;
        test_addr[1426] = 982;
        test_data[1426] = 33'd3325073124;
        test_addr[1427] = 983;
        test_data[1427] = 33'd253993433;
        test_addr[1428] = 984;
        test_data[1428] = 33'd1855044601;
        test_addr[1429] = 985;
        test_data[1429] = 33'd7299732777;
        test_addr[1430] = 986;
        test_data[1430] = 33'd4776303300;
        test_addr[1431] = 987;
        test_data[1431] = 33'd3846821607;
        test_addr[1432] = 988;
        test_data[1432] = 33'd6531544483;
        test_addr[1433] = 989;
        test_data[1433] = 33'd7170647933;
        test_addr[1434] = 990;
        test_data[1434] = 33'd76974876;
        test_addr[1435] = 991;
        test_data[1435] = 33'd7174531711;
        test_addr[1436] = 992;
        test_data[1436] = 33'd3935506262;
        test_addr[1437] = 993;
        test_data[1437] = 33'd4699311363;
        test_addr[1438] = 994;
        test_data[1438] = 33'd135589515;
        test_addr[1439] = 995;
        test_data[1439] = 33'd3833041508;
        test_addr[1440] = 996;
        test_data[1440] = 33'd744035756;
        test_addr[1441] = 997;
        test_data[1441] = 33'd6074174583;
        test_addr[1442] = 665;
        test_data[1442] = 33'd6063885606;
        test_addr[1443] = 666;
        test_data[1443] = 33'd1897257074;
        test_addr[1444] = 667;
        test_data[1444] = 33'd7173977800;
        test_addr[1445] = 668;
        test_data[1445] = 33'd3382879701;
        test_addr[1446] = 669;
        test_data[1446] = 33'd3165934849;
        test_addr[1447] = 670;
        test_data[1447] = 33'd2503869172;
        test_addr[1448] = 671;
        test_data[1448] = 33'd222714301;
        test_addr[1449] = 608;
        test_data[1449] = 33'd4136444716;
        test_addr[1450] = 609;
        test_data[1450] = 33'd8263265801;
        test_addr[1451] = 610;
        test_data[1451] = 33'd5076449630;
        test_addr[1452] = 611;
        test_data[1452] = 33'd2389840076;
        test_addr[1453] = 612;
        test_data[1453] = 33'd7927974040;
        test_addr[1454] = 613;
        test_data[1454] = 33'd2147567015;
        test_addr[1455] = 614;
        test_data[1455] = 33'd2943240457;
        test_addr[1456] = 615;
        test_data[1456] = 33'd4900340195;
        test_addr[1457] = 616;
        test_data[1457] = 33'd1345991342;
        test_addr[1458] = 617;
        test_data[1458] = 33'd979453922;
        test_addr[1459] = 618;
        test_data[1459] = 33'd7468868840;
        test_addr[1460] = 619;
        test_data[1460] = 33'd3667454584;
        test_addr[1461] = 620;
        test_data[1461] = 33'd2816982930;
        test_addr[1462] = 621;
        test_data[1462] = 33'd3470453698;
        test_addr[1463] = 622;
        test_data[1463] = 33'd3878932875;
        test_addr[1464] = 623;
        test_data[1464] = 33'd1284144988;
        test_addr[1465] = 624;
        test_data[1465] = 33'd7265078101;
        test_addr[1466] = 625;
        test_data[1466] = 33'd3243046981;
        test_addr[1467] = 626;
        test_data[1467] = 33'd2443222463;
        test_addr[1468] = 627;
        test_data[1468] = 33'd2341641585;
        test_addr[1469] = 628;
        test_data[1469] = 33'd4391894619;
        test_addr[1470] = 629;
        test_data[1470] = 33'd7253884188;
        test_addr[1471] = 630;
        test_data[1471] = 33'd2440170518;
        test_addr[1472] = 631;
        test_data[1472] = 33'd243801277;
        test_addr[1473] = 632;
        test_data[1473] = 33'd2564476576;
        test_addr[1474] = 633;
        test_data[1474] = 33'd916074034;
        test_addr[1475] = 634;
        test_data[1475] = 33'd3034116429;
        test_addr[1476] = 635;
        test_data[1476] = 33'd2142044604;
        test_addr[1477] = 636;
        test_data[1477] = 33'd3358336986;
        test_addr[1478] = 637;
        test_data[1478] = 33'd5107153102;
        test_addr[1479] = 672;
        test_data[1479] = 33'd336862564;
        test_addr[1480] = 673;
        test_data[1480] = 33'd4240157953;
        test_addr[1481] = 674;
        test_data[1481] = 33'd602961986;
        test_addr[1482] = 946;
        test_data[1482] = 33'd2617320100;
        test_addr[1483] = 947;
        test_data[1483] = 33'd1282791533;
        test_addr[1484] = 948;
        test_data[1484] = 33'd3621345128;
        test_addr[1485] = 949;
        test_data[1485] = 33'd3719719765;
        test_addr[1486] = 950;
        test_data[1486] = 33'd3002745736;
        test_addr[1487] = 951;
        test_data[1487] = 33'd52482036;
        test_addr[1488] = 675;
        test_data[1488] = 33'd953773948;
        test_addr[1489] = 676;
        test_data[1489] = 33'd7438577057;
        test_addr[1490] = 677;
        test_data[1490] = 33'd7807114274;
        test_addr[1491] = 100;
        test_data[1491] = 33'd8062810228;
        test_addr[1492] = 101;
        test_data[1492] = 33'd4476524971;
        test_addr[1493] = 102;
        test_data[1493] = 33'd4622918084;
        test_addr[1494] = 103;
        test_data[1494] = 33'd5451593796;
        test_addr[1495] = 678;
        test_data[1495] = 33'd2364391312;
        test_addr[1496] = 679;
        test_data[1496] = 33'd1418553768;
        test_addr[1497] = 680;
        test_data[1497] = 33'd6226246161;
        test_addr[1498] = 681;
        test_data[1498] = 33'd2488012861;
        test_addr[1499] = 682;
        test_data[1499] = 33'd7651004931;
        test_addr[1500] = 683;
        test_data[1500] = 33'd3868012904;
        test_addr[1501] = 684;
        test_data[1501] = 33'd878735113;
        test_addr[1502] = 685;
        test_data[1502] = 33'd1269636871;
        test_addr[1503] = 686;
        test_data[1503] = 33'd3201733946;
        test_addr[1504] = 687;
        test_data[1504] = 33'd1463662090;
        test_addr[1505] = 688;
        test_data[1505] = 33'd5879034205;
        test_addr[1506] = 689;
        test_data[1506] = 33'd743705583;
        test_addr[1507] = 690;
        test_data[1507] = 33'd2378395861;
        test_addr[1508] = 691;
        test_data[1508] = 33'd1508790809;
        test_addr[1509] = 692;
        test_data[1509] = 33'd735552833;
        test_addr[1510] = 693;
        test_data[1510] = 33'd6716960538;
        test_addr[1511] = 694;
        test_data[1511] = 33'd3269737490;
        test_addr[1512] = 695;
        test_data[1512] = 33'd6588594784;
        test_addr[1513] = 696;
        test_data[1513] = 33'd1822071661;
        test_addr[1514] = 697;
        test_data[1514] = 33'd1856755845;
        test_addr[1515] = 698;
        test_data[1515] = 33'd50727645;
        test_addr[1516] = 699;
        test_data[1516] = 33'd507075352;
        test_addr[1517] = 700;
        test_data[1517] = 33'd5076963731;
        test_addr[1518] = 701;
        test_data[1518] = 33'd2591022462;
        test_addr[1519] = 702;
        test_data[1519] = 33'd7664916829;
        test_addr[1520] = 703;
        test_data[1520] = 33'd2083865596;
        test_addr[1521] = 704;
        test_data[1521] = 33'd3483917983;
        test_addr[1522] = 705;
        test_data[1522] = 33'd6499083008;
        test_addr[1523] = 706;
        test_data[1523] = 33'd7107704823;
        test_addr[1524] = 707;
        test_data[1524] = 33'd7986234850;
        test_addr[1525] = 708;
        test_data[1525] = 33'd1052551570;
        test_addr[1526] = 709;
        test_data[1526] = 33'd3550218121;
        test_addr[1527] = 710;
        test_data[1527] = 33'd140022409;
        test_addr[1528] = 711;
        test_data[1528] = 33'd1464840222;
        test_addr[1529] = 712;
        test_data[1529] = 33'd5292868581;
        test_addr[1530] = 713;
        test_data[1530] = 33'd190684252;
        test_addr[1531] = 714;
        test_data[1531] = 33'd6688719563;
        test_addr[1532] = 715;
        test_data[1532] = 33'd4805767742;
        test_addr[1533] = 716;
        test_data[1533] = 33'd2485877949;
        test_addr[1534] = 717;
        test_data[1534] = 33'd5470387142;
        test_addr[1535] = 718;
        test_data[1535] = 33'd5043160793;
        test_addr[1536] = 552;
        test_data[1536] = 33'd5299066208;
        test_addr[1537] = 553;
        test_data[1537] = 33'd568073708;
        test_addr[1538] = 554;
        test_data[1538] = 33'd8250720715;
        test_addr[1539] = 555;
        test_data[1539] = 33'd8370111980;
        test_addr[1540] = 556;
        test_data[1540] = 33'd251347817;
        test_addr[1541] = 557;
        test_data[1541] = 33'd1317858012;
        test_addr[1542] = 558;
        test_data[1542] = 33'd7314714968;
        test_addr[1543] = 559;
        test_data[1543] = 33'd7352897182;
        test_addr[1544] = 560;
        test_data[1544] = 33'd7881743635;
        test_addr[1545] = 561;
        test_data[1545] = 33'd1077468732;
        test_addr[1546] = 562;
        test_data[1546] = 33'd579894608;
        test_addr[1547] = 719;
        test_data[1547] = 33'd3913089050;
        test_addr[1548] = 720;
        test_data[1548] = 33'd6783638668;
        test_addr[1549] = 721;
        test_data[1549] = 33'd6198622241;
        test_addr[1550] = 722;
        test_data[1550] = 33'd1996037175;
        test_addr[1551] = 723;
        test_data[1551] = 33'd485450652;
        test_addr[1552] = 737;
        test_data[1552] = 33'd3539109186;
        test_addr[1553] = 738;
        test_data[1553] = 33'd4807001843;
        test_addr[1554] = 739;
        test_data[1554] = 33'd3879861704;
        test_addr[1555] = 740;
        test_data[1555] = 33'd1695013347;
        test_addr[1556] = 741;
        test_data[1556] = 33'd7437458214;
        test_addr[1557] = 742;
        test_data[1557] = 33'd3001673332;
        test_addr[1558] = 724;
        test_data[1558] = 33'd3065873517;
        test_addr[1559] = 725;
        test_data[1559] = 33'd4231348663;
        test_addr[1560] = 726;
        test_data[1560] = 33'd4101723380;
        test_addr[1561] = 727;
        test_data[1561] = 33'd1097647790;
        test_addr[1562] = 728;
        test_data[1562] = 33'd3542905408;
        test_addr[1563] = 729;
        test_data[1563] = 33'd1951530555;
        test_addr[1564] = 730;
        test_data[1564] = 33'd5755265937;
        test_addr[1565] = 731;
        test_data[1565] = 33'd5268195625;
        test_addr[1566] = 732;
        test_data[1566] = 33'd1756047701;
        test_addr[1567] = 733;
        test_data[1567] = 33'd6586529010;
        test_addr[1568] = 734;
        test_data[1568] = 33'd5549199846;
        test_addr[1569] = 735;
        test_data[1569] = 33'd894928856;
        test_addr[1570] = 736;
        test_data[1570] = 33'd986423063;
        test_addr[1571] = 737;
        test_data[1571] = 33'd3539109186;
        test_addr[1572] = 738;
        test_data[1572] = 33'd512034547;
        test_addr[1573] = 185;
        test_data[1573] = 33'd4181767754;
        test_addr[1574] = 739;
        test_data[1574] = 33'd3879861704;
        test_addr[1575] = 740;
        test_data[1575] = 33'd1695013347;
        test_addr[1576] = 741;
        test_data[1576] = 33'd3142490918;
        test_addr[1577] = 742;
        test_data[1577] = 33'd3001673332;
        test_addr[1578] = 743;
        test_data[1578] = 33'd8198881353;
        test_addr[1579] = 744;
        test_data[1579] = 33'd1702935462;
        test_addr[1580] = 745;
        test_data[1580] = 33'd1433988871;
        test_addr[1581] = 746;
        test_data[1581] = 33'd3008884322;
        test_addr[1582] = 702;
        test_data[1582] = 33'd3369949533;
        test_addr[1583] = 747;
        test_data[1583] = 33'd740007894;
        test_addr[1584] = 748;
        test_data[1584] = 33'd6364794407;
        test_addr[1585] = 749;
        test_data[1585] = 33'd1788156813;
        test_addr[1586] = 750;
        test_data[1586] = 33'd80903859;
        test_addr[1587] = 751;
        test_data[1587] = 33'd2915964714;
        test_addr[1588] = 752;
        test_data[1588] = 33'd5281936767;
        test_addr[1589] = 753;
        test_data[1589] = 33'd2959231921;
        test_addr[1590] = 754;
        test_data[1590] = 33'd1522336256;
        test_addr[1591] = 755;
        test_data[1591] = 33'd6618786207;
        test_addr[1592] = 992;
        test_data[1592] = 33'd6352915573;
        test_addr[1593] = 993;
        test_data[1593] = 33'd5493523672;
        test_addr[1594] = 994;
        test_data[1594] = 33'd135589515;
        test_addr[1595] = 995;
        test_data[1595] = 33'd5497834178;
        test_addr[1596] = 996;
        test_data[1596] = 33'd744035756;
        test_addr[1597] = 997;
        test_data[1597] = 33'd1779207287;
        test_addr[1598] = 998;
        test_data[1598] = 33'd876875783;
        test_addr[1599] = 999;
        test_data[1599] = 33'd3854254352;
        test_addr[1600] = 756;
        test_data[1600] = 33'd4970434076;
        test_addr[1601] = 757;
        test_data[1601] = 33'd1411847050;
        test_addr[1602] = 758;
        test_data[1602] = 33'd8349285399;
        test_addr[1603] = 759;
        test_data[1603] = 33'd7022904326;
        test_addr[1604] = 760;
        test_data[1604] = 33'd5720971414;
        test_addr[1605] = 165;
        test_data[1605] = 33'd3249592251;
        test_addr[1606] = 166;
        test_data[1606] = 33'd1582126961;
        test_addr[1607] = 167;
        test_data[1607] = 33'd5075292357;
        test_addr[1608] = 168;
        test_data[1608] = 33'd3104257694;
        test_addr[1609] = 169;
        test_data[1609] = 33'd1157869169;
        test_addr[1610] = 170;
        test_data[1610] = 33'd983130549;
        test_addr[1611] = 171;
        test_data[1611] = 33'd5410923981;
        test_addr[1612] = 172;
        test_data[1612] = 33'd909425390;
        test_addr[1613] = 761;
        test_data[1613] = 33'd3442801664;
        test_addr[1614] = 526;
        test_data[1614] = 33'd324109075;
        test_addr[1615] = 527;
        test_data[1615] = 33'd3200519056;
        test_addr[1616] = 528;
        test_data[1616] = 33'd1322263514;
        test_addr[1617] = 529;
        test_data[1617] = 33'd1798434561;
        test_addr[1618] = 762;
        test_data[1618] = 33'd447989063;
        test_addr[1619] = 763;
        test_data[1619] = 33'd2202485930;
        test_addr[1620] = 764;
        test_data[1620] = 33'd2125336049;
        test_addr[1621] = 765;
        test_data[1621] = 33'd6666335522;
        test_addr[1622] = 766;
        test_data[1622] = 33'd2649969743;
        test_addr[1623] = 767;
        test_data[1623] = 33'd1956744276;
        test_addr[1624] = 768;
        test_data[1624] = 33'd5155258061;
        test_addr[1625] = 769;
        test_data[1625] = 33'd2812677734;
        test_addr[1626] = 770;
        test_data[1626] = 33'd4465541279;
        test_addr[1627] = 771;
        test_data[1627] = 33'd7314983127;
        test_addr[1628] = 772;
        test_data[1628] = 33'd1656105210;
        test_addr[1629] = 773;
        test_data[1629] = 33'd1846218975;
        test_addr[1630] = 774;
        test_data[1630] = 33'd3672349084;
        test_addr[1631] = 775;
        test_data[1631] = 33'd515219377;
        test_addr[1632] = 776;
        test_data[1632] = 33'd2726783519;
        test_addr[1633] = 543;
        test_data[1633] = 33'd6135567801;
        test_addr[1634] = 544;
        test_data[1634] = 33'd3366506315;
        test_addr[1635] = 545;
        test_data[1635] = 33'd2345963143;
        test_addr[1636] = 546;
        test_data[1636] = 33'd3228427618;
        test_addr[1637] = 777;
        test_data[1637] = 33'd6596750053;
        test_addr[1638] = 778;
        test_data[1638] = 33'd1166195020;
        test_addr[1639] = 779;
        test_data[1639] = 33'd2230018642;
        test_addr[1640] = 780;
        test_data[1640] = 33'd2527754555;
        test_addr[1641] = 781;
        test_data[1641] = 33'd6772934380;
        test_addr[1642] = 782;
        test_data[1642] = 33'd1898941484;
        test_addr[1643] = 783;
        test_data[1643] = 33'd8257152349;
        test_addr[1644] = 784;
        test_data[1644] = 33'd1886530748;
        test_addr[1645] = 785;
        test_data[1645] = 33'd1209496261;
        test_addr[1646] = 786;
        test_data[1646] = 33'd2215613352;
        test_addr[1647] = 787;
        test_data[1647] = 33'd8521166719;
        test_addr[1648] = 788;
        test_data[1648] = 33'd1647863726;
        test_addr[1649] = 789;
        test_data[1649] = 33'd1497512075;
        test_addr[1650] = 790;
        test_data[1650] = 33'd352952418;
        test_addr[1651] = 791;
        test_data[1651] = 33'd2708474774;
        test_addr[1652] = 792;
        test_data[1652] = 33'd2160729826;
        test_addr[1653] = 793;
        test_data[1653] = 33'd1811241968;
        test_addr[1654] = 794;
        test_data[1654] = 33'd3501008240;
        test_addr[1655] = 795;
        test_data[1655] = 33'd4091524596;
        test_addr[1656] = 796;
        test_data[1656] = 33'd1877609457;
        test_addr[1657] = 797;
        test_data[1657] = 33'd1827696675;
        test_addr[1658] = 798;
        test_data[1658] = 33'd3715808831;
        test_addr[1659] = 799;
        test_data[1659] = 33'd5366487588;
        test_addr[1660] = 800;
        test_data[1660] = 33'd356101764;
        test_addr[1661] = 801;
        test_data[1661] = 33'd4030133163;
        test_addr[1662] = 802;
        test_data[1662] = 33'd1172436856;
        test_addr[1663] = 803;
        test_data[1663] = 33'd3130885866;
        test_addr[1664] = 141;
        test_data[1664] = 33'd617480792;
        test_addr[1665] = 142;
        test_data[1665] = 33'd8030642561;
        test_addr[1666] = 143;
        test_data[1666] = 33'd3652162657;
        test_addr[1667] = 144;
        test_data[1667] = 33'd1695780936;
        test_addr[1668] = 145;
        test_data[1668] = 33'd3995848082;
        test_addr[1669] = 146;
        test_data[1669] = 33'd7480082207;
        test_addr[1670] = 804;
        test_data[1670] = 33'd1700099309;
        test_addr[1671] = 805;
        test_data[1671] = 33'd3103250482;
        test_addr[1672] = 806;
        test_data[1672] = 33'd2394794120;
        test_addr[1673] = 807;
        test_data[1673] = 33'd8058609481;
        test_addr[1674] = 808;
        test_data[1674] = 33'd8448028218;
        test_addr[1675] = 809;
        test_data[1675] = 33'd8235408708;
        test_addr[1676] = 810;
        test_data[1676] = 33'd1249729923;
        test_addr[1677] = 811;
        test_data[1677] = 33'd500276442;
        test_addr[1678] = 812;
        test_data[1678] = 33'd2198066108;
        test_addr[1679] = 813;
        test_data[1679] = 33'd1567399322;
        test_addr[1680] = 814;
        test_data[1680] = 33'd2725263772;
        test_addr[1681] = 815;
        test_data[1681] = 33'd1840551582;
        test_addr[1682] = 816;
        test_data[1682] = 33'd2266625000;
        test_addr[1683] = 817;
        test_data[1683] = 33'd6551114241;
        test_addr[1684] = 818;
        test_data[1684] = 33'd4127540968;
        test_addr[1685] = 819;
        test_data[1685] = 33'd7371068206;
        test_addr[1686] = 820;
        test_data[1686] = 33'd3540865897;
        test_addr[1687] = 821;
        test_data[1687] = 33'd2641923197;
        test_addr[1688] = 822;
        test_data[1688] = 33'd5615540270;
        test_addr[1689] = 823;
        test_data[1689] = 33'd803767947;
        test_addr[1690] = 824;
        test_data[1690] = 33'd3616832036;
        test_addr[1691] = 825;
        test_data[1691] = 33'd2843325391;
        test_addr[1692] = 826;
        test_data[1692] = 33'd1511462300;
        test_addr[1693] = 827;
        test_data[1693] = 33'd3433780831;
        test_addr[1694] = 828;
        test_data[1694] = 33'd3486781950;
        test_addr[1695] = 829;
        test_data[1695] = 33'd2744509025;
        test_addr[1696] = 830;
        test_data[1696] = 33'd2106790694;
        test_addr[1697] = 831;
        test_data[1697] = 33'd2989084624;
        test_addr[1698] = 832;
        test_data[1698] = 33'd636608990;
        test_addr[1699] = 833;
        test_data[1699] = 33'd2060550887;
        test_addr[1700] = 834;
        test_data[1700] = 33'd2565041108;
        test_addr[1701] = 835;
        test_data[1701] = 33'd2346246843;
        test_addr[1702] = 580;
        test_data[1702] = 33'd7015096091;
        test_addr[1703] = 581;
        test_data[1703] = 33'd2909404543;
        test_addr[1704] = 582;
        test_data[1704] = 33'd7467296719;
        test_addr[1705] = 583;
        test_data[1705] = 33'd7531187025;
        test_addr[1706] = 836;
        test_data[1706] = 33'd374999801;
        test_addr[1707] = 837;
        test_data[1707] = 33'd2883404476;
        test_addr[1708] = 838;
        test_data[1708] = 33'd1505196816;
        test_addr[1709] = 839;
        test_data[1709] = 33'd5737299357;
        test_addr[1710] = 840;
        test_data[1710] = 33'd1961400636;
        test_addr[1711] = 841;
        test_data[1711] = 33'd6372796827;
        test_addr[1712] = 842;
        test_data[1712] = 33'd8588963328;
        test_addr[1713] = 843;
        test_data[1713] = 33'd6304832363;
        test_addr[1714] = 844;
        test_data[1714] = 33'd3760661512;
        test_addr[1715] = 623;
        test_data[1715] = 33'd1284144988;
        test_addr[1716] = 624;
        test_data[1716] = 33'd2970110805;
        test_addr[1717] = 625;
        test_data[1717] = 33'd3243046981;
        test_addr[1718] = 626;
        test_data[1718] = 33'd2443222463;
        test_addr[1719] = 845;
        test_data[1719] = 33'd2007080822;
        test_addr[1720] = 846;
        test_data[1720] = 33'd2513345585;
        test_addr[1721] = 847;
        test_data[1721] = 33'd8150960161;
        test_addr[1722] = 848;
        test_data[1722] = 33'd4157002771;
        test_addr[1723] = 849;
        test_data[1723] = 33'd1713558479;
        test_addr[1724] = 774;
        test_data[1724] = 33'd3672349084;
        test_addr[1725] = 775;
        test_data[1725] = 33'd515219377;
        test_addr[1726] = 776;
        test_data[1726] = 33'd6171296466;
        test_addr[1727] = 777;
        test_data[1727] = 33'd2301782757;
        test_addr[1728] = 778;
        test_data[1728] = 33'd1166195020;
        test_addr[1729] = 779;
        test_data[1729] = 33'd2230018642;
        test_addr[1730] = 780;
        test_data[1730] = 33'd2527754555;
        test_addr[1731] = 781;
        test_data[1731] = 33'd2477967084;
        test_addr[1732] = 782;
        test_data[1732] = 33'd1898941484;
        test_addr[1733] = 783;
        test_data[1733] = 33'd3962185053;
        test_addr[1734] = 784;
        test_data[1734] = 33'd1886530748;
        test_addr[1735] = 785;
        test_data[1735] = 33'd6387051819;
        test_addr[1736] = 786;
        test_data[1736] = 33'd8129373253;
        test_addr[1737] = 787;
        test_data[1737] = 33'd4226199423;
        test_addr[1738] = 788;
        test_data[1738] = 33'd1647863726;
        test_addr[1739] = 789;
        test_data[1739] = 33'd1497512075;
        test_addr[1740] = 790;
        test_data[1740] = 33'd7156766762;
        test_addr[1741] = 791;
        test_data[1741] = 33'd2708474774;
        test_addr[1742] = 792;
        test_data[1742] = 33'd2160729826;
        test_addr[1743] = 793;
        test_data[1743] = 33'd8092136419;
        test_addr[1744] = 794;
        test_data[1744] = 33'd3501008240;
        test_addr[1745] = 795;
        test_data[1745] = 33'd7593209422;
        test_addr[1746] = 796;
        test_data[1746] = 33'd8040900152;
        test_addr[1747] = 797;
        test_data[1747] = 33'd7395010893;
        test_addr[1748] = 798;
        test_data[1748] = 33'd3715808831;
        test_addr[1749] = 799;
        test_data[1749] = 33'd8469407695;
        test_addr[1750] = 800;
        test_data[1750] = 33'd356101764;
        test_addr[1751] = 801;
        test_data[1751] = 33'd4030133163;
        test_addr[1752] = 802;
        test_data[1752] = 33'd6290786249;
        test_addr[1753] = 803;
        test_data[1753] = 33'd3130885866;
        test_addr[1754] = 804;
        test_data[1754] = 33'd7738768642;
        test_addr[1755] = 805;
        test_data[1755] = 33'd8268326549;
        test_addr[1756] = 850;
        test_data[1756] = 33'd8316028576;
        test_addr[1757] = 851;
        test_data[1757] = 33'd5272172544;
        test_addr[1758] = 852;
        test_data[1758] = 33'd309025837;
        test_addr[1759] = 853;
        test_data[1759] = 33'd7836171202;
        test_addr[1760] = 854;
        test_data[1760] = 33'd6932907730;
        test_addr[1761] = 855;
        test_data[1761] = 33'd3556722367;
        test_addr[1762] = 856;
        test_data[1762] = 33'd4744016863;
        test_addr[1763] = 857;
        test_data[1763] = 33'd5231986222;
        test_addr[1764] = 858;
        test_data[1764] = 33'd5450132936;
        test_addr[1765] = 859;
        test_data[1765] = 33'd61833049;
        test_addr[1766] = 860;
        test_data[1766] = 33'd542097023;
        test_addr[1767] = 861;
        test_data[1767] = 33'd4331106816;
        test_addr[1768] = 862;
        test_data[1768] = 33'd6831312161;
        test_addr[1769] = 863;
        test_data[1769] = 33'd1939476593;
        test_addr[1770] = 864;
        test_data[1770] = 33'd7973984885;
        test_addr[1771] = 865;
        test_data[1771] = 33'd2384212187;
        test_addr[1772] = 866;
        test_data[1772] = 33'd6362850299;
        test_addr[1773] = 867;
        test_data[1773] = 33'd5699323080;
        test_addr[1774] = 868;
        test_data[1774] = 33'd3122240770;
        test_addr[1775] = 869;
        test_data[1775] = 33'd7684597002;
        test_addr[1776] = 870;
        test_data[1776] = 33'd2534380821;
        test_addr[1777] = 871;
        test_data[1777] = 33'd6678578740;
        test_addr[1778] = 371;
        test_data[1778] = 33'd338135865;
        test_addr[1779] = 372;
        test_data[1779] = 33'd605321337;
        test_addr[1780] = 373;
        test_data[1780] = 33'd1524839362;
        test_addr[1781] = 374;
        test_data[1781] = 33'd3597032391;
        test_addr[1782] = 375;
        test_data[1782] = 33'd86563587;
        test_addr[1783] = 376;
        test_data[1783] = 33'd2007598323;
        test_addr[1784] = 377;
        test_data[1784] = 33'd7787542567;
        test_addr[1785] = 378;
        test_data[1785] = 33'd1683535556;
        test_addr[1786] = 379;
        test_data[1786] = 33'd6367333343;
        test_addr[1787] = 380;
        test_data[1787] = 33'd931778438;
        test_addr[1788] = 381;
        test_data[1788] = 33'd5443954104;
        test_addr[1789] = 382;
        test_data[1789] = 33'd3335835945;
        test_addr[1790] = 383;
        test_data[1790] = 33'd51573383;
        test_addr[1791] = 384;
        test_data[1791] = 33'd5704310455;
        test_addr[1792] = 385;
        test_data[1792] = 33'd2749730789;
        test_addr[1793] = 386;
        test_data[1793] = 33'd8253538334;
        test_addr[1794] = 387;
        test_data[1794] = 33'd1682531476;
        test_addr[1795] = 872;
        test_data[1795] = 33'd1325586264;
        test_addr[1796] = 873;
        test_data[1796] = 33'd2396752366;
        test_addr[1797] = 199;
        test_data[1797] = 33'd7149632812;
        test_addr[1798] = 874;
        test_data[1798] = 33'd25727163;
        test_addr[1799] = 875;
        test_data[1799] = 33'd477340108;
        test_addr[1800] = 876;
        test_data[1800] = 33'd6118708650;
        test_addr[1801] = 877;
        test_data[1801] = 33'd3703124324;
        test_addr[1802] = 878;
        test_data[1802] = 33'd7455681220;
        test_addr[1803] = 879;
        test_data[1803] = 33'd1464330775;
        test_addr[1804] = 880;
        test_data[1804] = 33'd5125152461;
        test_addr[1805] = 881;
        test_data[1805] = 33'd1506016935;
        test_addr[1806] = 882;
        test_data[1806] = 33'd3835130572;
        test_addr[1807] = 883;
        test_data[1807] = 33'd3004317571;
        test_addr[1808] = 884;
        test_data[1808] = 33'd422576570;
        test_addr[1809] = 885;
        test_data[1809] = 33'd7137560792;
        test_addr[1810] = 886;
        test_data[1810] = 33'd4672651606;
        test_addr[1811] = 887;
        test_data[1811] = 33'd3092087050;
        test_addr[1812] = 888;
        test_data[1812] = 33'd309666434;
        test_addr[1813] = 889;
        test_data[1813] = 33'd955985398;
        test_addr[1814] = 890;
        test_data[1814] = 33'd3259517725;
        test_addr[1815] = 891;
        test_data[1815] = 33'd514451412;
        test_addr[1816] = 892;
        test_data[1816] = 33'd1499118016;
        test_addr[1817] = 893;
        test_data[1817] = 33'd2707802790;
        test_addr[1818] = 894;
        test_data[1818] = 33'd5533347990;
        test_addr[1819] = 895;
        test_data[1819] = 33'd653469184;
        test_addr[1820] = 896;
        test_data[1820] = 33'd1456229272;
        test_addr[1821] = 897;
        test_data[1821] = 33'd7171973589;
        test_addr[1822] = 898;
        test_data[1822] = 33'd1668711176;
        test_addr[1823] = 899;
        test_data[1823] = 33'd7714134038;
        test_addr[1824] = 900;
        test_data[1824] = 33'd2401073967;
        test_addr[1825] = 901;
        test_data[1825] = 33'd3853423062;
        test_addr[1826] = 902;
        test_data[1826] = 33'd3321083730;
        test_addr[1827] = 903;
        test_data[1827] = 33'd3146695517;
        test_addr[1828] = 904;
        test_data[1828] = 33'd2772309859;
        test_addr[1829] = 905;
        test_data[1829] = 33'd6696899773;
        test_addr[1830] = 906;
        test_data[1830] = 33'd3531140847;
        test_addr[1831] = 907;
        test_data[1831] = 33'd1045330292;
        test_addr[1832] = 908;
        test_data[1832] = 33'd6490352387;
        test_addr[1833] = 909;
        test_data[1833] = 33'd1069087929;
        test_addr[1834] = 910;
        test_data[1834] = 33'd3676552037;
        test_addr[1835] = 911;
        test_data[1835] = 33'd284526649;
        test_addr[1836] = 912;
        test_data[1836] = 33'd1888499141;
        test_addr[1837] = 913;
        test_data[1837] = 33'd714474144;
        test_addr[1838] = 914;
        test_data[1838] = 33'd1975795592;
        test_addr[1839] = 915;
        test_data[1839] = 33'd4165669295;
        test_addr[1840] = 916;
        test_data[1840] = 33'd6189185498;
        test_addr[1841] = 917;
        test_data[1841] = 33'd6723366678;
        test_addr[1842] = 918;
        test_data[1842] = 33'd4239968030;
        test_addr[1843] = 919;
        test_data[1843] = 33'd2730893660;
        test_addr[1844] = 920;
        test_data[1844] = 33'd3606140741;
        test_addr[1845] = 921;
        test_data[1845] = 33'd662140256;
        test_addr[1846] = 922;
        test_data[1846] = 33'd6560833774;
        test_addr[1847] = 923;
        test_data[1847] = 33'd1827564675;
        test_addr[1848] = 924;
        test_data[1848] = 33'd6504497535;
        test_addr[1849] = 925;
        test_data[1849] = 33'd164526863;
        test_addr[1850] = 926;
        test_data[1850] = 33'd2588329358;
        test_addr[1851] = 927;
        test_data[1851] = 33'd2111508981;
        test_addr[1852] = 928;
        test_data[1852] = 33'd6845141849;
        test_addr[1853] = 929;
        test_data[1853] = 33'd4115151129;
        test_addr[1854] = 930;
        test_data[1854] = 33'd3058555497;
        test_addr[1855] = 931;
        test_data[1855] = 33'd7928129;
        test_addr[1856] = 932;
        test_data[1856] = 33'd1498951355;
        test_addr[1857] = 933;
        test_data[1857] = 33'd4583631697;
        test_addr[1858] = 934;
        test_data[1858] = 33'd3936725344;
        test_addr[1859] = 935;
        test_data[1859] = 33'd3119130326;
        test_addr[1860] = 936;
        test_data[1860] = 33'd6224241231;
        test_addr[1861] = 937;
        test_data[1861] = 33'd4402459234;
        test_addr[1862] = 938;
        test_data[1862] = 33'd3703155137;
        test_addr[1863] = 939;
        test_data[1863] = 33'd889180094;
        test_addr[1864] = 940;
        test_data[1864] = 33'd7146597005;
        test_addr[1865] = 941;
        test_data[1865] = 33'd1981406870;
        test_addr[1866] = 942;
        test_data[1866] = 33'd2606351839;
        test_addr[1867] = 943;
        test_data[1867] = 33'd3360306346;
        test_addr[1868] = 944;
        test_data[1868] = 33'd134171436;
        test_addr[1869] = 945;
        test_data[1869] = 33'd3068243404;
        test_addr[1870] = 946;
        test_data[1870] = 33'd2617320100;
        test_addr[1871] = 947;
        test_data[1871] = 33'd1282791533;
        test_addr[1872] = 948;
        test_data[1872] = 33'd4380437515;
        test_addr[1873] = 949;
        test_data[1873] = 33'd7542680554;
        test_addr[1874] = 950;
        test_data[1874] = 33'd8211421438;
        test_addr[1875] = 951;
        test_data[1875] = 33'd4618431132;
        test_addr[1876] = 952;
        test_data[1876] = 33'd3444183392;
        test_addr[1877] = 993;
        test_data[1877] = 33'd1198556376;
        test_addr[1878] = 994;
        test_data[1878] = 33'd135589515;
        test_addr[1879] = 995;
        test_data[1879] = 33'd6925513095;
        test_addr[1880] = 996;
        test_data[1880] = 33'd4565465161;
        test_addr[1881] = 997;
        test_data[1881] = 33'd1779207287;
        test_addr[1882] = 998;
        test_data[1882] = 33'd876875783;
        test_addr[1883] = 999;
        test_data[1883] = 33'd3854254352;
        test_addr[1884] = 1000;
        test_data[1884] = 33'd3694084155;
        test_addr[1885] = 1001;
        test_data[1885] = 33'd249958146;
        test_addr[1886] = 1002;
        test_data[1886] = 33'd6705521369;
        test_addr[1887] = 953;
        test_data[1887] = 33'd702849432;
        test_addr[1888] = 954;
        test_data[1888] = 33'd247955198;
        test_addr[1889] = 955;
        test_data[1889] = 33'd6012998518;
        test_addr[1890] = 956;
        test_data[1890] = 33'd5967415152;
        test_addr[1891] = 957;
        test_data[1891] = 33'd2402321614;
        test_addr[1892] = 516;
        test_data[1892] = 33'd5294562905;
        test_addr[1893] = 517;
        test_data[1893] = 33'd162263759;
        test_addr[1894] = 518;
        test_data[1894] = 33'd48984368;
        test_addr[1895] = 519;
        test_data[1895] = 33'd1574109177;
        test_addr[1896] = 520;
        test_data[1896] = 33'd847712690;
        test_addr[1897] = 521;
        test_data[1897] = 33'd7282052445;
        test_addr[1898] = 522;
        test_data[1898] = 33'd6788729351;
        test_addr[1899] = 523;
        test_data[1899] = 33'd40985424;
        test_addr[1900] = 524;
        test_data[1900] = 33'd3607396520;
        test_addr[1901] = 525;
        test_data[1901] = 33'd3236712843;
        test_addr[1902] = 526;
        test_data[1902] = 33'd7178597925;
        test_addr[1903] = 527;
        test_data[1903] = 33'd4951700111;
        test_addr[1904] = 528;
        test_data[1904] = 33'd8270216597;
        test_addr[1905] = 529;
        test_data[1905] = 33'd6794523113;
        test_addr[1906] = 958;
        test_data[1906] = 33'd3879054770;
        test_addr[1907] = 959;
        test_data[1907] = 33'd4485440417;
        test_addr[1908] = 960;
        test_data[1908] = 33'd6208656204;
        test_addr[1909] = 961;
        test_data[1909] = 33'd7732740071;
        test_addr[1910] = 962;
        test_data[1910] = 33'd4548740606;
        test_addr[1911] = 963;
        test_data[1911] = 33'd5323410519;
        test_addr[1912] = 964;
        test_data[1912] = 33'd881417507;
        test_addr[1913] = 965;
        test_data[1913] = 33'd8356678199;
        test_addr[1914] = 966;
        test_data[1914] = 33'd3326283328;
        test_addr[1915] = 967;
        test_data[1915] = 33'd2283602290;
        test_addr[1916] = 968;
        test_data[1916] = 33'd380593856;
        test_addr[1917] = 969;
        test_data[1917] = 33'd2228588555;
        test_addr[1918] = 970;
        test_data[1918] = 33'd5483164390;
        test_addr[1919] = 971;
        test_data[1919] = 33'd2956302870;
        test_addr[1920] = 972;
        test_data[1920] = 33'd1407407298;
        test_addr[1921] = 973;
        test_data[1921] = 33'd214877909;
        test_addr[1922] = 974;
        test_data[1922] = 33'd1727455379;
        test_addr[1923] = 975;
        test_data[1923] = 33'd3749386507;
        test_addr[1924] = 976;
        test_data[1924] = 33'd7862093385;
        test_addr[1925] = 977;
        test_data[1925] = 33'd892255078;
        test_addr[1926] = 978;
        test_data[1926] = 33'd2804270651;
        test_addr[1927] = 979;
        test_data[1927] = 33'd3376760179;
        test_addr[1928] = 980;
        test_data[1928] = 33'd8021453663;
        test_addr[1929] = 981;
        test_data[1929] = 33'd4566466225;
        test_addr[1930] = 982;
        test_data[1930] = 33'd8319695347;
        test_addr[1931] = 983;
        test_data[1931] = 33'd253993433;
        test_addr[1932] = 984;
        test_data[1932] = 33'd7505752309;
        test_addr[1933] = 166;
        test_data[1933] = 33'd5448102248;
        test_addr[1934] = 985;
        test_data[1934] = 33'd3004765481;
        test_addr[1935] = 986;
        test_data[1935] = 33'd481336004;
        test_addr[1936] = 987;
        test_data[1936] = 33'd3846821607;
        test_addr[1937] = 988;
        test_data[1937] = 33'd2236577187;
        test_addr[1938] = 308;
        test_data[1938] = 33'd8567279930;
        test_addr[1939] = 309;
        test_data[1939] = 33'd7331472381;
        test_addr[1940] = 310;
        test_data[1940] = 33'd892285550;
        test_addr[1941] = 311;
        test_data[1941] = 33'd757719279;
        test_addr[1942] = 312;
        test_data[1942] = 33'd1581510545;
        test_addr[1943] = 313;
        test_data[1943] = 33'd5370165080;
        test_addr[1944] = 314;
        test_data[1944] = 33'd7736352701;
        test_addr[1945] = 315;
        test_data[1945] = 33'd1538426196;
        test_addr[1946] = 316;
        test_data[1946] = 33'd2469986364;
        test_addr[1947] = 317;
        test_data[1947] = 33'd5702258048;
        test_addr[1948] = 318;
        test_data[1948] = 33'd3064576727;
        test_addr[1949] = 319;
        test_data[1949] = 33'd8197986863;
        test_addr[1950] = 320;
        test_data[1950] = 33'd8055818287;
        test_addr[1951] = 321;
        test_data[1951] = 33'd2227829365;
        test_addr[1952] = 322;
        test_data[1952] = 33'd2533921378;
        test_addr[1953] = 323;
        test_data[1953] = 33'd5918440114;
        test_addr[1954] = 324;
        test_data[1954] = 33'd2565321190;
        test_addr[1955] = 325;
        test_data[1955] = 33'd2573803079;
        test_addr[1956] = 326;
        test_data[1956] = 33'd8209596303;
        test_addr[1957] = 327;
        test_data[1957] = 33'd2931519176;
        test_addr[1958] = 328;
        test_data[1958] = 33'd6673572259;
        test_addr[1959] = 329;
        test_data[1959] = 33'd3283575319;
        test_addr[1960] = 330;
        test_data[1960] = 33'd3377953911;
        test_addr[1961] = 331;
        test_data[1961] = 33'd4985951395;
        test_addr[1962] = 332;
        test_data[1962] = 33'd403124710;
        test_addr[1963] = 333;
        test_data[1963] = 33'd7239578651;
        test_addr[1964] = 334;
        test_data[1964] = 33'd2841628197;
        test_addr[1965] = 335;
        test_data[1965] = 33'd4393672975;
        test_addr[1966] = 336;
        test_data[1966] = 33'd745322449;
        test_addr[1967] = 337;
        test_data[1967] = 33'd4218420959;
        test_addr[1968] = 338;
        test_data[1968] = 33'd2832891657;
        test_addr[1969] = 339;
        test_data[1969] = 33'd3237287086;
        test_addr[1970] = 340;
        test_data[1970] = 33'd2309224711;
        test_addr[1971] = 989;
        test_data[1971] = 33'd2875680637;
        test_addr[1972] = 990;
        test_data[1972] = 33'd76974876;
        test_addr[1973] = 991;
        test_data[1973] = 33'd2879564415;
        test_addr[1974] = 961;
        test_data[1974] = 33'd3437772775;
        test_addr[1975] = 962;
        test_data[1975] = 33'd8423752763;
        test_addr[1976] = 963;
        test_data[1976] = 33'd1028443223;
        test_addr[1977] = 964;
        test_data[1977] = 33'd881417507;
        test_addr[1978] = 992;
        test_data[1978] = 33'd5003295842;
        test_addr[1979] = 993;
        test_data[1979] = 33'd1198556376;
        test_addr[1980] = 994;
        test_data[1980] = 33'd135589515;
        test_addr[1981] = 995;
        test_data[1981] = 33'd2630545799;
        test_addr[1982] = 996;
        test_data[1982] = 33'd6543041539;
        test_addr[1983] = 583;
        test_data[1983] = 33'd7586922318;
        test_addr[1984] = 584;
        test_data[1984] = 33'd602235759;
        test_addr[1985] = 997;
        test_data[1985] = 33'd1779207287;
        test_addr[1986] = 998;
        test_data[1986] = 33'd876875783;
        test_addr[1987] = 119;
        test_data[1987] = 33'd2347492591;
        test_addr[1988] = 120;
        test_data[1988] = 33'd5910634323;
        test_addr[1989] = 121;
        test_data[1989] = 33'd1116625760;
        test_addr[1990] = 122;
        test_data[1990] = 33'd2382385405;
        test_addr[1991] = 123;
        test_data[1991] = 33'd2378157637;
        test_addr[1992] = 124;
        test_data[1992] = 33'd1884814149;
        test_addr[1993] = 125;
        test_data[1993] = 33'd2085264057;
        test_addr[1994] = 126;
        test_data[1994] = 33'd5639093396;
        test_addr[1995] = 127;
        test_data[1995] = 33'd7385180007;
        test_addr[1996] = 128;
        test_data[1996] = 33'd8342257270;
        test_addr[1997] = 129;
        test_data[1997] = 33'd2800001925;
        test_addr[1998] = 130;
        test_data[1998] = 33'd1440556275;
        test_addr[1999] = 131;
        test_data[1999] = 33'd3900854079;
        test_addr[2000] = 132;
        test_data[2000] = 33'd1523580593;
        test_addr[2001] = 133;
        test_data[2001] = 33'd2214113554;
        test_addr[2002] = 134;
        test_data[2002] = 33'd137763915;
        test_addr[2003] = 135;
        test_data[2003] = 33'd1350958361;
        test_addr[2004] = 136;
        test_data[2004] = 33'd7253872385;
        test_addr[2005] = 137;
        test_data[2005] = 33'd2021339031;
        test_addr[2006] = 138;
        test_data[2006] = 33'd7220872979;
        test_addr[2007] = 139;
        test_data[2007] = 33'd5067202422;
        test_addr[2008] = 140;
        test_data[2008] = 33'd6303628706;
        test_addr[2009] = 141;
        test_data[2009] = 33'd4825128796;
        test_addr[2010] = 999;
        test_data[2010] = 33'd3854254352;
        test_addr[2011] = 1000;
        test_data[2011] = 33'd6402717314;
        test_addr[2012] = 1001;
        test_data[2012] = 33'd7043951130;
        test_addr[2013] = 1002;
        test_data[2013] = 33'd5623543198;
        test_addr[2014] = 1003;
        test_data[2014] = 33'd4769314635;
        test_addr[2015] = 1004;
        test_data[2015] = 33'd7173304410;
        test_addr[2016] = 1005;
        test_data[2016] = 33'd7702450674;
        test_addr[2017] = 1006;
        test_data[2017] = 33'd6253881499;
        test_addr[2018] = 1007;
        test_data[2018] = 33'd7326211608;
        test_addr[2019] = 1008;
        test_data[2019] = 33'd2879552693;
        test_addr[2020] = 1009;
        test_data[2020] = 33'd4292225377;
        test_addr[2021] = 1010;
        test_data[2021] = 33'd3905914762;
        test_addr[2022] = 504;
        test_data[2022] = 33'd1574083226;
        test_addr[2023] = 505;
        test_data[2023] = 33'd7321205044;
        test_addr[2024] = 506;
        test_data[2024] = 33'd4602611477;
        test_addr[2025] = 507;
        test_data[2025] = 33'd7012156211;
        test_addr[2026] = 508;
        test_data[2026] = 33'd3420814826;
        test_addr[2027] = 509;
        test_data[2027] = 33'd282828349;
        test_addr[2028] = 1011;
        test_data[2028] = 33'd4682166737;
        test_addr[2029] = 1012;
        test_data[2029] = 33'd6892099853;
        test_addr[2030] = 992;
        test_data[2030] = 33'd708328546;
        test_addr[2031] = 993;
        test_data[2031] = 33'd8104316790;
        test_addr[2032] = 994;
        test_data[2032] = 33'd135589515;
        test_addr[2033] = 995;
        test_data[2033] = 33'd2630545799;
        test_addr[2034] = 996;
        test_data[2034] = 33'd2248074243;
        test_addr[2035] = 997;
        test_data[2035] = 33'd1779207287;
        test_addr[2036] = 998;
        test_data[2036] = 33'd876875783;
        test_addr[2037] = 999;
        test_data[2037] = 33'd3854254352;
        test_addr[2038] = 1000;
        test_data[2038] = 33'd8511935471;
        test_addr[2039] = 1001;
        test_data[2039] = 33'd2748983834;
        test_addr[2040] = 1002;
        test_data[2040] = 33'd1328575902;
        test_addr[2041] = 1003;
        test_data[2041] = 33'd6769463651;
        test_addr[2042] = 1004;
        test_data[2042] = 33'd2878337114;
        test_addr[2043] = 1005;
        test_data[2043] = 33'd3407483378;
        test_addr[2044] = 1006;
        test_data[2044] = 33'd1958914203;
        test_addr[2045] = 1007;
        test_data[2045] = 33'd5591189562;
        test_addr[2046] = 1013;
        test_data[2046] = 33'd2767383358;
        test_addr[2047] = 41;
        test_data[2047] = 33'd897063482;
        test_addr[2048] = 42;
        test_data[2048] = 33'd6613643249;
        test_addr[2049] = 43;
        test_data[2049] = 33'd2262236211;
        test_addr[2050] = 44;
        test_data[2050] = 33'd5873660969;
        test_addr[2051] = 45;
        test_data[2051] = 33'd3465150654;
        test_addr[2052] = 46;
        test_data[2052] = 33'd3718565962;
        test_addr[2053] = 47;
        test_data[2053] = 33'd456343954;
        test_addr[2054] = 48;
        test_data[2054] = 33'd6905215262;
        test_addr[2055] = 49;
        test_data[2055] = 33'd6269774836;
        test_addr[2056] = 50;
        test_data[2056] = 33'd6248446704;
        test_addr[2057] = 51;
        test_data[2057] = 33'd7156242608;
        test_addr[2058] = 52;
        test_data[2058] = 33'd6379180833;
        test_addr[2059] = 53;
        test_data[2059] = 33'd1099507616;
        test_addr[2060] = 54;
        test_data[2060] = 33'd5781160086;
        test_addr[2061] = 55;
        test_data[2061] = 33'd855085249;
        test_addr[2062] = 56;
        test_data[2062] = 33'd7497968234;
        test_addr[2063] = 57;
        test_data[2063] = 33'd3178846984;
        test_addr[2064] = 58;
        test_data[2064] = 33'd8271984641;
        test_addr[2065] = 59;
        test_data[2065] = 33'd3097027422;
        test_addr[2066] = 60;
        test_data[2066] = 33'd8370575873;
        test_addr[2067] = 1014;
        test_data[2067] = 33'd2467778259;
        test_addr[2068] = 56;
        test_data[2068] = 33'd3203000938;
        test_addr[2069] = 57;
        test_data[2069] = 33'd4981033431;
        test_addr[2070] = 58;
        test_data[2070] = 33'd3977017345;
        test_addr[2071] = 1015;
        test_data[2071] = 33'd1385438272;
        test_addr[2072] = 1016;
        test_data[2072] = 33'd659905488;
        test_addr[2073] = 1017;
        test_data[2073] = 33'd4843047852;
        test_addr[2074] = 1018;
        test_data[2074] = 33'd1719465706;
        test_addr[2075] = 1019;
        test_data[2075] = 33'd4716771183;
        test_addr[2076] = 1020;
        test_data[2076] = 33'd1493206180;
        test_addr[2077] = 1021;
        test_data[2077] = 33'd349429309;
        test_addr[2078] = 1022;
        test_data[2078] = 33'd2782636993;
        test_addr[2079] = 1023;
        test_data[2079] = 33'd1545197175;
        test_addr[2080] = 0;
        test_data[2080] = 33'd1052567479;
        test_addr[2081] = 1;
        test_data[2081] = 33'd3962591981;
        test_addr[2082] = 2;
        test_data[2082] = 33'd4750023242;
        test_addr[2083] = 3;
        test_data[2083] = 33'd3048570618;
        test_addr[2084] = 4;
        test_data[2084] = 33'd2553106968;
        test_addr[2085] = 5;
        test_data[2085] = 33'd5342572551;
        test_addr[2086] = 6;
        test_data[2086] = 33'd4900443055;
        test_addr[2087] = 7;
        test_data[2087] = 33'd3045195451;
        test_addr[2088] = 8;
        test_data[2088] = 33'd606447009;
        test_addr[2089] = 9;
        test_data[2089] = 33'd5532300043;
        test_addr[2090] = 10;
        test_data[2090] = 33'd93493361;
        test_addr[2091] = 11;
        test_data[2091] = 33'd4541805971;
        test_addr[2092] = 12;
        test_data[2092] = 33'd770777372;
        test_addr[2093] = 13;
        test_data[2093] = 33'd675467997;
        test_addr[2094] = 14;
        test_data[2094] = 33'd1785532064;
        test_addr[2095] = 15;
        test_data[2095] = 33'd1461300596;
        test_addr[2096] = 700;
        test_data[2096] = 33'd781996435;
        test_addr[2097] = 701;
        test_data[2097] = 33'd2591022462;
        test_addr[2098] = 702;
        test_data[2098] = 33'd6684205556;
        test_addr[2099] = 703;
        test_data[2099] = 33'd2083865596;
        test_addr[2100] = 16;
        test_data[2100] = 33'd1426394555;
        test_addr[2101] = 17;
        test_data[2101] = 33'd5486861288;
        test_addr[2102] = 18;
        test_data[2102] = 33'd3721935424;
        test_addr[2103] = 19;
        test_data[2103] = 33'd5435458901;
        test_addr[2104] = 20;
        test_data[2104] = 33'd6117406119;
        test_addr[2105] = 21;
        test_data[2105] = 33'd1976287339;
        test_addr[2106] = 22;
        test_data[2106] = 33'd7139625494;
        test_addr[2107] = 23;
        test_data[2107] = 33'd6117860919;
        test_addr[2108] = 24;
        test_data[2108] = 33'd6288025823;
        test_addr[2109] = 25;
        test_data[2109] = 33'd5234388798;
        test_addr[2110] = 26;
        test_data[2110] = 33'd59093393;
        test_addr[2111] = 97;
        test_data[2111] = 33'd8563907445;
        test_addr[2112] = 98;
        test_data[2112] = 33'd2187286926;
        test_addr[2113] = 27;
        test_data[2113] = 33'd1793516677;
        test_addr[2114] = 28;
        test_data[2114] = 33'd3711284261;
        test_addr[2115] = 436;
        test_data[2115] = 33'd4273322909;
        test_addr[2116] = 437;
        test_data[2116] = 33'd1332405155;
        test_addr[2117] = 438;
        test_data[2117] = 33'd2165787536;
        test_addr[2118] = 439;
        test_data[2118] = 33'd1956260871;
        test_addr[2119] = 440;
        test_data[2119] = 33'd7332949487;
        test_addr[2120] = 441;
        test_data[2120] = 33'd65904936;
        test_addr[2121] = 442;
        test_data[2121] = 33'd8465290642;
        test_addr[2122] = 443;
        test_data[2122] = 33'd1076063113;
        test_addr[2123] = 444;
        test_data[2123] = 33'd4084632541;
        test_addr[2124] = 445;
        test_data[2124] = 33'd6022292004;
        test_addr[2125] = 446;
        test_data[2125] = 33'd2468389652;
        test_addr[2126] = 447;
        test_data[2126] = 33'd7671614534;
        test_addr[2127] = 448;
        test_data[2127] = 33'd1265298441;
        test_addr[2128] = 449;
        test_data[2128] = 33'd2908833870;
        test_addr[2129] = 450;
        test_data[2129] = 33'd2162667854;
        test_addr[2130] = 29;
        test_data[2130] = 33'd3303147092;
        test_addr[2131] = 30;
        test_data[2131] = 33'd6433108521;
        test_addr[2132] = 31;
        test_data[2132] = 33'd1352203701;
        test_addr[2133] = 106;
        test_data[2133] = 33'd7603460943;
        test_addr[2134] = 107;
        test_data[2134] = 33'd2778245487;
        test_addr[2135] = 108;
        test_data[2135] = 33'd2932393469;
        test_addr[2136] = 109;
        test_data[2136] = 33'd664815512;
        test_addr[2137] = 32;
        test_data[2137] = 33'd6856416775;
        test_addr[2138] = 33;
        test_data[2138] = 33'd3582404842;
        test_addr[2139] = 34;
        test_data[2139] = 33'd3140383792;
        test_addr[2140] = 74;
        test_data[2140] = 33'd2454510322;
        test_addr[2141] = 75;
        test_data[2141] = 33'd1791303464;
        test_addr[2142] = 76;
        test_data[2142] = 33'd3925384761;
        test_addr[2143] = 77;
        test_data[2143] = 33'd3109637631;
        test_addr[2144] = 78;
        test_data[2144] = 33'd728046435;
        test_addr[2145] = 79;
        test_data[2145] = 33'd3563875528;
        test_addr[2146] = 80;
        test_data[2146] = 33'd3205303345;
        test_addr[2147] = 81;
        test_data[2147] = 33'd7100122818;
        test_addr[2148] = 82;
        test_data[2148] = 33'd4356747263;
        test_addr[2149] = 35;
        test_data[2149] = 33'd1823217833;
        test_addr[2150] = 36;
        test_data[2150] = 33'd7993197846;
        test_addr[2151] = 37;
        test_data[2151] = 33'd1883382384;
        test_addr[2152] = 38;
        test_data[2152] = 33'd982384382;
        test_addr[2153] = 39;
        test_data[2153] = 33'd5457644941;
        test_addr[2154] = 40;
        test_data[2154] = 33'd334310572;
        test_addr[2155] = 41;
        test_data[2155] = 33'd897063482;
        test_addr[2156] = 42;
        test_data[2156] = 33'd4967229546;
        test_addr[2157] = 43;
        test_data[2157] = 33'd2262236211;
        test_addr[2158] = 491;
        test_data[2158] = 33'd2354554954;
        test_addr[2159] = 492;
        test_data[2159] = 33'd2825740953;
        test_addr[2160] = 493;
        test_data[2160] = 33'd5203967599;
        test_addr[2161] = 494;
        test_data[2161] = 33'd5457069258;
        test_addr[2162] = 495;
        test_data[2162] = 33'd7320772597;
        test_addr[2163] = 496;
        test_data[2163] = 33'd7312378447;
        test_addr[2164] = 44;
        test_data[2164] = 33'd1578693673;
        test_addr[2165] = 994;
        test_data[2165] = 33'd6646876598;
        test_addr[2166] = 995;
        test_data[2166] = 33'd6284517811;
        test_addr[2167] = 996;
        test_data[2167] = 33'd2248074243;
        test_addr[2168] = 997;
        test_data[2168] = 33'd4515373366;
        test_addr[2169] = 998;
        test_data[2169] = 33'd5773394048;
        test_addr[2170] = 999;
        test_data[2170] = 33'd3854254352;
        test_addr[2171] = 1000;
        test_data[2171] = 33'd5592614810;
        test_addr[2172] = 1001;
        test_data[2172] = 33'd2748983834;
        test_addr[2173] = 1002;
        test_data[2173] = 33'd1328575902;
        test_addr[2174] = 1003;
        test_data[2174] = 33'd2474496355;
        test_addr[2175] = 1004;
        test_data[2175] = 33'd5079463595;
        test_addr[2176] = 1005;
        test_data[2176] = 33'd3407483378;
        test_addr[2177] = 1006;
        test_data[2177] = 33'd1958914203;
        test_addr[2178] = 1007;
        test_data[2178] = 33'd8079719326;
        test_addr[2179] = 1008;
        test_data[2179] = 33'd4752287400;
        test_addr[2180] = 1009;
        test_data[2180] = 33'd7792233376;
        test_addr[2181] = 1010;
        test_data[2181] = 33'd3905914762;
        test_addr[2182] = 1011;
        test_data[2182] = 33'd7079457773;
        test_addr[2183] = 1012;
        test_data[2183] = 33'd6934339880;
        test_addr[2184] = 1013;
        test_data[2184] = 33'd4742756179;
        test_addr[2185] = 1014;
        test_data[2185] = 33'd2467778259;
        test_addr[2186] = 1015;
        test_data[2186] = 33'd1385438272;
        test_addr[2187] = 1016;
        test_data[2187] = 33'd5640454915;
        test_addr[2188] = 45;
        test_data[2188] = 33'd3465150654;
        test_addr[2189] = 46;
        test_data[2189] = 33'd3718565962;
        test_addr[2190] = 47;
        test_data[2190] = 33'd5403954007;
        test_addr[2191] = 48;
        test_data[2191] = 33'd2610247966;
        test_addr[2192] = 49;
        test_data[2192] = 33'd4748157793;
        test_addr[2193] = 50;
        test_data[2193] = 33'd4599731446;
        test_addr[2194] = 51;
        test_data[2194] = 33'd2861275312;
        test_addr[2195] = 52;
        test_data[2195] = 33'd2084213537;
        test_addr[2196] = 53;
        test_data[2196] = 33'd5261437822;
        test_addr[2197] = 54;
        test_data[2197] = 33'd4550810783;
        test_addr[2198] = 55;
        test_data[2198] = 33'd5073567813;
        test_addr[2199] = 56;
        test_data[2199] = 33'd6835015880;
        test_addr[2200] = 57;
        test_data[2200] = 33'd686066135;
        test_addr[2201] = 58;
        test_data[2201] = 33'd6738921515;
        test_addr[2202] = 59;
        test_data[2202] = 33'd5045232051;
        test_addr[2203] = 60;
        test_data[2203] = 33'd4075608577;
        test_addr[2204] = 61;
        test_data[2204] = 33'd468031354;
        test_addr[2205] = 62;
        test_data[2205] = 33'd209881339;
        test_addr[2206] = 63;
        test_data[2206] = 33'd4681755784;
        test_addr[2207] = 64;
        test_data[2207] = 33'd819283579;
        test_addr[2208] = 65;
        test_data[2208] = 33'd3395724500;
        test_addr[2209] = 66;
        test_data[2209] = 33'd2714239827;
        test_addr[2210] = 67;
        test_data[2210] = 33'd5486797767;
        test_addr[2211] = 68;
        test_data[2211] = 33'd5487790991;
        test_addr[2212] = 69;
        test_data[2212] = 33'd2018933038;
        test_addr[2213] = 170;
        test_data[2213] = 33'd6989569287;
        test_addr[2214] = 171;
        test_data[2214] = 33'd1115956685;
        test_addr[2215] = 172;
        test_data[2215] = 33'd909425390;
        test_addr[2216] = 173;
        test_data[2216] = 33'd3560746765;
        test_addr[2217] = 174;
        test_data[2217] = 33'd6698560639;
        test_addr[2218] = 70;
        test_data[2218] = 33'd1396858963;
        test_addr[2219] = 71;
        test_data[2219] = 33'd3173125001;
        test_addr[2220] = 72;
        test_data[2220] = 33'd5751546395;
        test_addr[2221] = 73;
        test_data[2221] = 33'd546788671;
        test_addr[2222] = 74;
        test_data[2222] = 33'd2454510322;
        test_addr[2223] = 75;
        test_data[2223] = 33'd1791303464;
        test_addr[2224] = 76;
        test_data[2224] = 33'd3925384761;
        test_addr[2225] = 77;
        test_data[2225] = 33'd3109637631;
        test_addr[2226] = 78;
        test_data[2226] = 33'd728046435;
        test_addr[2227] = 79;
        test_data[2227] = 33'd3563875528;
        test_addr[2228] = 80;
        test_data[2228] = 33'd4325539926;
        test_addr[2229] = 117;
        test_data[2229] = 33'd2384278837;
        test_addr[2230] = 118;
        test_data[2230] = 33'd6459911056;
        test_addr[2231] = 81;
        test_data[2231] = 33'd2805155522;
        test_addr[2232] = 82;
        test_data[2232] = 33'd61779967;
        test_addr[2233] = 83;
        test_data[2233] = 33'd1065113936;
        test_addr[2234] = 84;
        test_data[2234] = 33'd6395548261;
        test_addr[2235] = 85;
        test_data[2235] = 33'd3558159285;
        test_addr[2236] = 86;
        test_data[2236] = 33'd3378272531;
        test_addr[2237] = 87;
        test_data[2237] = 33'd2963060552;
        test_addr[2238] = 88;
        test_data[2238] = 33'd8003817043;
        test_addr[2239] = 89;
        test_data[2239] = 33'd8002085915;
        test_addr[2240] = 90;
        test_data[2240] = 33'd7707031542;
        test_addr[2241] = 91;
        test_data[2241] = 33'd7243474396;
        test_addr[2242] = 92;
        test_data[2242] = 33'd242469961;
        test_addr[2243] = 93;
        test_data[2243] = 33'd93622177;
        test_addr[2244] = 94;
        test_data[2244] = 33'd8388456601;
        test_addr[2245] = 95;
        test_data[2245] = 33'd4186162648;
        test_addr[2246] = 96;
        test_data[2246] = 33'd1514847775;
        test_addr[2247] = 97;
        test_data[2247] = 33'd6200325465;
        test_addr[2248] = 98;
        test_data[2248] = 33'd2187286926;
        test_addr[2249] = 470;
        test_data[2249] = 33'd1434334882;
        test_addr[2250] = 471;
        test_data[2250] = 33'd5291622033;
        test_addr[2251] = 472;
        test_data[2251] = 33'd173483137;
        test_addr[2252] = 473;
        test_data[2252] = 33'd3858581669;
        test_addr[2253] = 474;
        test_data[2253] = 33'd242718291;
        test_addr[2254] = 99;
        test_data[2254] = 33'd3901445798;
        test_addr[2255] = 100;
        test_data[2255] = 33'd3767842932;
        test_addr[2256] = 101;
        test_data[2256] = 33'd181557675;
        test_addr[2257] = 102;
        test_data[2257] = 33'd6910263211;
        test_addr[2258] = 889;
        test_data[2258] = 33'd6388966396;
        test_addr[2259] = 890;
        test_data[2259] = 33'd6169865098;
        test_addr[2260] = 891;
        test_data[2260] = 33'd514451412;
        test_addr[2261] = 892;
        test_data[2261] = 33'd1499118016;
        test_addr[2262] = 893;
        test_data[2262] = 33'd2707802790;
        test_addr[2263] = 894;
        test_data[2263] = 33'd5303623324;
        test_addr[2264] = 895;
        test_data[2264] = 33'd653469184;
        test_addr[2265] = 896;
        test_data[2265] = 33'd7684930131;
        test_addr[2266] = 897;
        test_data[2266] = 33'd5079532296;
        test_addr[2267] = 898;
        test_data[2267] = 33'd1668711176;
        test_addr[2268] = 899;
        test_data[2268] = 33'd3419166742;
        test_addr[2269] = 900;
        test_data[2269] = 33'd2401073967;
        test_addr[2270] = 901;
        test_data[2270] = 33'd6725991954;
        test_addr[2271] = 902;
        test_data[2271] = 33'd5410072963;
        test_addr[2272] = 903;
        test_data[2272] = 33'd3146695517;
        test_addr[2273] = 904;
        test_data[2273] = 33'd2772309859;
        test_addr[2274] = 905;
        test_data[2274] = 33'd2401932477;
        test_addr[2275] = 103;
        test_data[2275] = 33'd1156626500;
        test_addr[2276] = 104;
        test_data[2276] = 33'd2137822137;
        test_addr[2277] = 105;
        test_data[2277] = 33'd7757510027;
        test_addr[2278] = 106;
        test_data[2278] = 33'd7529718783;
        test_addr[2279] = 107;
        test_data[2279] = 33'd6940015076;
        test_addr[2280] = 108;
        test_data[2280] = 33'd2932393469;
        test_addr[2281] = 109;
        test_data[2281] = 33'd664815512;
        test_addr[2282] = 110;
        test_data[2282] = 33'd8201328566;
        test_addr[2283] = 395;
        test_data[2283] = 33'd101142806;
        test_addr[2284] = 396;
        test_data[2284] = 33'd3707484179;
        test_addr[2285] = 111;
        test_data[2285] = 33'd2870920926;
        test_addr[2286] = 112;
        test_data[2286] = 33'd53516149;
        test_addr[2287] = 113;
        test_data[2287] = 33'd6501103629;
        test_addr[2288] = 114;
        test_data[2288] = 33'd574419132;
        test_addr[2289] = 115;
        test_data[2289] = 33'd4921273943;
        test_addr[2290] = 116;
        test_data[2290] = 33'd7877370868;
        test_addr[2291] = 117;
        test_data[2291] = 33'd2384278837;
        test_addr[2292] = 118;
        test_data[2292] = 33'd2164943760;
        test_addr[2293] = 119;
        test_data[2293] = 33'd8099199264;
        test_addr[2294] = 120;
        test_data[2294] = 33'd5141250520;
        test_addr[2295] = 121;
        test_data[2295] = 33'd5578495447;
        test_addr[2296] = 122;
        test_data[2296] = 33'd2382385405;
        test_addr[2297] = 123;
        test_data[2297] = 33'd7490057119;
        test_addr[2298] = 124;
        test_data[2298] = 33'd1884814149;
        test_addr[2299] = 125;
        test_data[2299] = 33'd2085264057;
        test_addr[2300] = 126;
        test_data[2300] = 33'd1344126100;
        test_addr[2301] = 127;
        test_data[2301] = 33'd3090212711;
        test_addr[2302] = 128;
        test_data[2302] = 33'd7707224920;
        test_addr[2303] = 129;
        test_data[2303] = 33'd5838542161;
        test_addr[2304] = 130;
        test_data[2304] = 33'd8338297321;
        test_addr[2305] = 131;
        test_data[2305] = 33'd3900854079;
        test_addr[2306] = 132;
        test_data[2306] = 33'd1523580593;
        test_addr[2307] = 133;
        test_data[2307] = 33'd5419534436;
        test_addr[2308] = 134;
        test_data[2308] = 33'd137763915;
        test_addr[2309] = 135;
        test_data[2309] = 33'd7080602654;
        test_addr[2310] = 136;
        test_data[2310] = 33'd2958905089;
        test_addr[2311] = 137;
        test_data[2311] = 33'd2021339031;
        test_addr[2312] = 138;
        test_data[2312] = 33'd2925905683;
        test_addr[2313] = 139;
        test_data[2313] = 33'd772235126;
        test_addr[2314] = 140;
        test_data[2314] = 33'd5934557254;
        test_addr[2315] = 474;
        test_data[2315] = 33'd8116031455;
        test_addr[2316] = 475;
        test_data[2316] = 33'd3328634438;
        test_addr[2317] = 476;
        test_data[2317] = 33'd2866816344;
        test_addr[2318] = 477;
        test_data[2318] = 33'd3782855187;
        test_addr[2319] = 478;
        test_data[2319] = 33'd7358705249;
        test_addr[2320] = 479;
        test_data[2320] = 33'd2293417793;
        test_addr[2321] = 480;
        test_data[2321] = 33'd799026300;
        test_addr[2322] = 481;
        test_data[2322] = 33'd3611509395;
        test_addr[2323] = 482;
        test_data[2323] = 33'd107901289;
        test_addr[2324] = 483;
        test_data[2324] = 33'd7067809590;
        test_addr[2325] = 484;
        test_data[2325] = 33'd8331985314;
        test_addr[2326] = 485;
        test_data[2326] = 33'd453359906;
        test_addr[2327] = 486;
        test_data[2327] = 33'd4650647886;
        test_addr[2328] = 487;
        test_data[2328] = 33'd3658540064;
        test_addr[2329] = 488;
        test_data[2329] = 33'd6847399823;
        test_addr[2330] = 141;
        test_data[2330] = 33'd530161500;
        test_addr[2331] = 142;
        test_data[2331] = 33'd7945804192;
        test_addr[2332] = 143;
        test_data[2332] = 33'd3652162657;
        test_addr[2333] = 144;
        test_data[2333] = 33'd1695780936;
        test_addr[2334] = 752;
        test_data[2334] = 33'd4524138811;
        test_addr[2335] = 145;
        test_data[2335] = 33'd3995848082;
        test_addr[2336] = 146;
        test_data[2336] = 33'd5684245726;
        test_addr[2337] = 147;
        test_data[2337] = 33'd776585138;
        test_addr[2338] = 148;
        test_data[2338] = 33'd1157076026;
        test_addr[2339] = 149;
        test_data[2339] = 33'd4440064177;
        test_addr[2340] = 150;
        test_data[2340] = 33'd6263918358;
        test_addr[2341] = 151;
        test_data[2341] = 33'd8320134126;
        test_addr[2342] = 152;
        test_data[2342] = 33'd5612302050;
        test_addr[2343] = 153;
        test_data[2343] = 33'd3554490906;
        test_addr[2344] = 154;
        test_data[2344] = 33'd3756857754;
        test_addr[2345] = 155;
        test_data[2345] = 33'd2556299901;
        test_addr[2346] = 156;
        test_data[2346] = 33'd6867276875;
        test_addr[2347] = 157;
        test_data[2347] = 33'd7151779014;
        test_addr[2348] = 158;
        test_data[2348] = 33'd5431168201;
        test_addr[2349] = 159;
        test_data[2349] = 33'd8292200285;
        test_addr[2350] = 160;
        test_data[2350] = 33'd688845184;
        test_addr[2351] = 578;
        test_data[2351] = 33'd2578797357;
        test_addr[2352] = 579;
        test_data[2352] = 33'd6879461314;
        test_addr[2353] = 580;
        test_data[2353] = 33'd2720128795;
        test_addr[2354] = 581;
        test_data[2354] = 33'd2909404543;
        test_addr[2355] = 582;
        test_data[2355] = 33'd3172329423;
        test_addr[2356] = 583;
        test_data[2356] = 33'd5809302311;
        test_addr[2357] = 584;
        test_data[2357] = 33'd6789904915;
        test_addr[2358] = 585;
        test_data[2358] = 33'd3545634013;
        test_addr[2359] = 586;
        test_data[2359] = 33'd3351735354;
        test_addr[2360] = 587;
        test_data[2360] = 33'd291280601;
        test_addr[2361] = 588;
        test_data[2361] = 33'd2023990209;
        test_addr[2362] = 589;
        test_data[2362] = 33'd8551072231;
        test_addr[2363] = 161;
        test_data[2363] = 33'd1723706081;
        test_addr[2364] = 162;
        test_data[2364] = 33'd5906723659;
        test_addr[2365] = 163;
        test_data[2365] = 33'd3158758932;
        test_addr[2366] = 164;
        test_data[2366] = 33'd10763549;
        test_addr[2367] = 165;
        test_data[2367] = 33'd3249592251;
        test_addr[2368] = 166;
        test_data[2368] = 33'd1153134952;
        test_addr[2369] = 167;
        test_data[2369] = 33'd780325061;
        test_addr[2370] = 168;
        test_data[2370] = 33'd5287624587;
        test_addr[2371] = 169;
        test_data[2371] = 33'd1157869169;
        test_addr[2372] = 170;
        test_data[2372] = 33'd8346260430;
        test_addr[2373] = 171;
        test_data[2373] = 33'd1115956685;
        test_addr[2374] = 172;
        test_data[2374] = 33'd7166282654;
        test_addr[2375] = 173;
        test_data[2375] = 33'd3560746765;
        test_addr[2376] = 174;
        test_data[2376] = 33'd5378616378;
        test_addr[2377] = 419;
        test_data[2377] = 33'd3137721503;
        test_addr[2378] = 420;
        test_data[2378] = 33'd1115528034;
        test_addr[2379] = 421;
        test_data[2379] = 33'd749396176;
        test_addr[2380] = 422;
        test_data[2380] = 33'd4129404128;
        test_addr[2381] = 423;
        test_data[2381] = 33'd6631864797;
        test_addr[2382] = 424;
        test_data[2382] = 33'd4259167484;
        test_addr[2383] = 425;
        test_data[2383] = 33'd7727562116;
        test_addr[2384] = 426;
        test_data[2384] = 33'd7782393828;
        test_addr[2385] = 175;
        test_data[2385] = 33'd5196918124;
        test_addr[2386] = 176;
        test_data[2386] = 33'd1240149642;
        test_addr[2387] = 177;
        test_data[2387] = 33'd1530014160;
        test_addr[2388] = 178;
        test_data[2388] = 33'd3395508098;
        test_addr[2389] = 179;
        test_data[2389] = 33'd2165023982;
        test_addr[2390] = 180;
        test_data[2390] = 33'd54599123;
        test_addr[2391] = 181;
        test_data[2391] = 33'd7857480347;
        test_addr[2392] = 182;
        test_data[2392] = 33'd830768617;
        test_addr[2393] = 183;
        test_data[2393] = 33'd818267281;
        test_addr[2394] = 184;
        test_data[2394] = 33'd2586566993;
        test_addr[2395] = 874;
        test_data[2395] = 33'd25727163;
        test_addr[2396] = 875;
        test_data[2396] = 33'd477340108;
        test_addr[2397] = 876;
        test_data[2397] = 33'd1823741354;
        test_addr[2398] = 877;
        test_data[2398] = 33'd3703124324;
        test_addr[2399] = 878;
        test_data[2399] = 33'd3160713924;
        test_addr[2400] = 879;
        test_data[2400] = 33'd1464330775;
        test_addr[2401] = 185;
        test_data[2401] = 33'd4181767754;
        test_addr[2402] = 186;
        test_data[2402] = 33'd3269096103;
        test_addr[2403] = 187;
        test_data[2403] = 33'd640249350;
        test_addr[2404] = 188;
        test_data[2404] = 33'd3301553819;
        test_addr[2405] = 189;
        test_data[2405] = 33'd966409649;
        test_addr[2406] = 190;
        test_data[2406] = 33'd1159409871;
        test_addr[2407] = 191;
        test_data[2407] = 33'd3743401526;
        test_addr[2408] = 192;
        test_data[2408] = 33'd1686812042;
        test_addr[2409] = 193;
        test_data[2409] = 33'd389818431;
        test_addr[2410] = 194;
        test_data[2410] = 33'd6790167650;
        test_addr[2411] = 195;
        test_data[2411] = 33'd6033207716;
        test_addr[2412] = 504;
        test_data[2412] = 33'd1574083226;
        test_addr[2413] = 196;
        test_data[2413] = 33'd871728998;
        test_addr[2414] = 197;
        test_data[2414] = 33'd3233146207;
        test_addr[2415] = 198;
        test_data[2415] = 33'd1825329058;
        test_addr[2416] = 199;
        test_data[2416] = 33'd2854665516;
        test_addr[2417] = 200;
        test_data[2417] = 33'd4473735638;
        test_addr[2418] = 201;
        test_data[2418] = 33'd3380527101;
        test_addr[2419] = 202;
        test_data[2419] = 33'd1247379816;
        test_addr[2420] = 203;
        test_data[2420] = 33'd6425686896;
        test_addr[2421] = 204;
        test_data[2421] = 33'd1243827460;
        test_addr[2422] = 205;
        test_data[2422] = 33'd2438118847;
        test_addr[2423] = 206;
        test_data[2423] = 33'd5795108548;
        test_addr[2424] = 207;
        test_data[2424] = 33'd867306624;
        test_addr[2425] = 208;
        test_data[2425] = 33'd738706595;
        test_addr[2426] = 209;
        test_data[2426] = 33'd4188964105;
        test_addr[2427] = 210;
        test_data[2427] = 33'd7234543531;
        test_addr[2428] = 211;
        test_data[2428] = 33'd1230764576;
        test_addr[2429] = 212;
        test_data[2429] = 33'd3427452440;
        test_addr[2430] = 213;
        test_data[2430] = 33'd4895730682;
        test_addr[2431] = 214;
        test_data[2431] = 33'd8470526789;
        test_addr[2432] = 215;
        test_data[2432] = 33'd8523703255;
        test_addr[2433] = 216;
        test_data[2433] = 33'd6269712273;
        test_addr[2434] = 217;
        test_data[2434] = 33'd91812431;
        test_addr[2435] = 218;
        test_data[2435] = 33'd709857341;
        test_addr[2436] = 219;
        test_data[2436] = 33'd2099384420;
        test_addr[2437] = 220;
        test_data[2437] = 33'd3956104701;
        test_addr[2438] = 221;
        test_data[2438] = 33'd2513170581;
        test_addr[2439] = 222;
        test_data[2439] = 33'd8249509419;
        test_addr[2440] = 223;
        test_data[2440] = 33'd1645865683;
        test_addr[2441] = 224;
        test_data[2441] = 33'd4306876234;
        test_addr[2442] = 225;
        test_data[2442] = 33'd1888744485;
        test_addr[2443] = 226;
        test_data[2443] = 33'd8368298845;
        test_addr[2444] = 227;
        test_data[2444] = 33'd7331059257;
        test_addr[2445] = 228;
        test_data[2445] = 33'd6088129208;
        test_addr[2446] = 229;
        test_data[2446] = 33'd1524904068;
        test_addr[2447] = 230;
        test_data[2447] = 33'd5924708617;
        test_addr[2448] = 231;
        test_data[2448] = 33'd3982051426;
        test_addr[2449] = 232;
        test_data[2449] = 33'd274384184;
        test_addr[2450] = 233;
        test_data[2450] = 33'd312253816;
        test_addr[2451] = 234;
        test_data[2451] = 33'd8351468584;
        test_addr[2452] = 815;
        test_data[2452] = 33'd1840551582;
        test_addr[2453] = 816;
        test_data[2453] = 33'd2266625000;
        test_addr[2454] = 817;
        test_data[2454] = 33'd2256146945;
        test_addr[2455] = 818;
        test_data[2455] = 33'd4127540968;
        test_addr[2456] = 819;
        test_data[2456] = 33'd3076100910;
        test_addr[2457] = 820;
        test_data[2457] = 33'd5018783740;
        test_addr[2458] = 821;
        test_data[2458] = 33'd2641923197;
        test_addr[2459] = 822;
        test_data[2459] = 33'd1320572974;
        test_addr[2460] = 235;
        test_data[2460] = 33'd2756285415;
        test_addr[2461] = 236;
        test_data[2461] = 33'd2037725383;
        test_addr[2462] = 237;
        test_data[2462] = 33'd1838823857;
        test_addr[2463] = 238;
        test_data[2463] = 33'd3263906087;
        test_addr[2464] = 239;
        test_data[2464] = 33'd5230782008;
        test_addr[2465] = 240;
        test_data[2465] = 33'd5838189927;
        test_addr[2466] = 241;
        test_data[2466] = 33'd3949767492;
        test_addr[2467] = 242;
        test_data[2467] = 33'd136386603;
        test_addr[2468] = 243;
        test_data[2468] = 33'd8173554433;
        test_addr[2469] = 244;
        test_data[2469] = 33'd7776842285;
        test_addr[2470] = 245;
        test_data[2470] = 33'd1169530796;
        test_addr[2471] = 246;
        test_data[2471] = 33'd4612705530;
        test_addr[2472] = 247;
        test_data[2472] = 33'd4279741554;
        test_addr[2473] = 980;
        test_data[2473] = 33'd7343423938;
        test_addr[2474] = 981;
        test_data[2474] = 33'd271498929;
        test_addr[2475] = 982;
        test_data[2475] = 33'd4024728051;
        test_addr[2476] = 983;
        test_data[2476] = 33'd253993433;
        test_addr[2477] = 984;
        test_data[2477] = 33'd6559262834;
        test_addr[2478] = 985;
        test_data[2478] = 33'd3004765481;
        test_addr[2479] = 986;
        test_data[2479] = 33'd481336004;
        test_addr[2480] = 987;
        test_data[2480] = 33'd5037197853;
        test_addr[2481] = 988;
        test_data[2481] = 33'd2236577187;
        test_addr[2482] = 989;
        test_data[2482] = 33'd5305087530;
        test_addr[2483] = 990;
        test_data[2483] = 33'd76974876;
        test_addr[2484] = 991;
        test_data[2484] = 33'd2879564415;
        test_addr[2485] = 992;
        test_data[2485] = 33'd708328546;
        test_addr[2486] = 993;
        test_data[2486] = 33'd3809349494;
        test_addr[2487] = 994;
        test_data[2487] = 33'd2351909302;
        test_addr[2488] = 995;
        test_data[2488] = 33'd1989550515;
        test_addr[2489] = 996;
        test_data[2489] = 33'd2248074243;
        test_addr[2490] = 997;
        test_data[2490] = 33'd220406070;
        test_addr[2491] = 998;
        test_data[2491] = 33'd1478426752;
        test_addr[2492] = 999;
        test_data[2492] = 33'd6898264891;
        test_addr[2493] = 1000;
        test_data[2493] = 33'd1297647514;
        test_addr[2494] = 1001;
        test_data[2494] = 33'd2748983834;
        test_addr[2495] = 248;
        test_data[2495] = 33'd3051279083;
        test_addr[2496] = 249;
        test_data[2496] = 33'd8433309260;
        test_addr[2497] = 250;
        test_data[2497] = 33'd7279977767;
        test_addr[2498] = 251;
        test_data[2498] = 33'd3980764503;
        test_addr[2499] = 252;
        test_data[2499] = 33'd2162877397;
        test_addr[2500] = 253;
        test_data[2500] = 33'd3083274420;
        test_addr[2501] = 254;
        test_data[2501] = 33'd7813357341;
        test_addr[2502] = 255;
        test_data[2502] = 33'd3333567760;
        test_addr[2503] = 256;
        test_data[2503] = 33'd5980419491;
        test_addr[2504] = 257;
        test_data[2504] = 33'd6853674203;
        test_addr[2505] = 258;
        test_data[2505] = 33'd4966550398;
        test_addr[2506] = 259;
        test_data[2506] = 33'd5667705617;
        test_addr[2507] = 260;
        test_data[2507] = 33'd3517079168;
        test_addr[2508] = 261;
        test_data[2508] = 33'd1946819819;
        test_addr[2509] = 262;
        test_data[2509] = 33'd6227461944;
        test_addr[2510] = 263;
        test_data[2510] = 33'd997948274;
        test_addr[2511] = 264;
        test_data[2511] = 33'd247406431;
        test_addr[2512] = 265;
        test_data[2512] = 33'd4016900671;
        test_addr[2513] = 266;
        test_data[2513] = 33'd1955864689;
        test_addr[2514] = 267;
        test_data[2514] = 33'd2384171014;
        test_addr[2515] = 268;
        test_data[2515] = 33'd4135890016;
        test_addr[2516] = 269;
        test_data[2516] = 33'd1870362431;
        test_addr[2517] = 270;
        test_data[2517] = 33'd3591863440;
        test_addr[2518] = 271;
        test_data[2518] = 33'd4531310315;
        test_addr[2519] = 272;
        test_data[2519] = 33'd1532962167;
        test_addr[2520] = 273;
        test_data[2520] = 33'd1672741610;
        test_addr[2521] = 51;
        test_data[2521] = 33'd2861275312;
        test_addr[2522] = 52;
        test_data[2522] = 33'd2084213537;
        test_addr[2523] = 274;
        test_data[2523] = 33'd2078674897;
        test_addr[2524] = 275;
        test_data[2524] = 33'd2726176411;
        test_addr[2525] = 276;
        test_data[2525] = 33'd2588319835;
        test_addr[2526] = 277;
        test_data[2526] = 33'd7563975946;
        test_addr[2527] = 278;
        test_data[2527] = 33'd976419527;
        test_addr[2528] = 279;
        test_data[2528] = 33'd3323213134;
        test_addr[2529] = 280;
        test_data[2529] = 33'd6066536715;
        test_addr[2530] = 281;
        test_data[2530] = 33'd5081925649;
        test_addr[2531] = 282;
        test_data[2531] = 33'd643220710;
        test_addr[2532] = 283;
        test_data[2532] = 33'd1833786499;
        test_addr[2533] = 284;
        test_data[2533] = 33'd1308087725;
        test_addr[2534] = 285;
        test_data[2534] = 33'd554349352;
        test_addr[2535] = 286;
        test_data[2535] = 33'd5491165863;
        test_addr[2536] = 287;
        test_data[2536] = 33'd3928208796;
        test_addr[2537] = 288;
        test_data[2537] = 33'd1952811514;
        test_addr[2538] = 289;
        test_data[2538] = 33'd3503208650;
        test_addr[2539] = 290;
        test_data[2539] = 33'd8118036607;
        test_addr[2540] = 291;
        test_data[2540] = 33'd5564642805;
        test_addr[2541] = 292;
        test_data[2541] = 33'd7604449387;
        test_addr[2542] = 293;
        test_data[2542] = 33'd8335756129;
        test_addr[2543] = 294;
        test_data[2543] = 33'd1462825451;
        test_addr[2544] = 295;
        test_data[2544] = 33'd6192801395;
        test_addr[2545] = 296;
        test_data[2545] = 33'd1858975900;
        test_addr[2546] = 297;
        test_data[2546] = 33'd1255568382;
        test_addr[2547] = 298;
        test_data[2547] = 33'd1354822540;
        test_addr[2548] = 299;
        test_data[2548] = 33'd6584826213;
        test_addr[2549] = 300;
        test_data[2549] = 33'd8479837476;
        test_addr[2550] = 301;
        test_data[2550] = 33'd7631830210;
        test_addr[2551] = 302;
        test_data[2551] = 33'd5528476766;
        test_addr[2552] = 303;
        test_data[2552] = 33'd7725836185;
        test_addr[2553] = 304;
        test_data[2553] = 33'd3131755163;
        test_addr[2554] = 305;
        test_data[2554] = 33'd2985268612;
        test_addr[2555] = 306;
        test_data[2555] = 33'd2048220064;
        test_addr[2556] = 307;
        test_data[2556] = 33'd395268976;
        test_addr[2557] = 308;
        test_data[2557] = 33'd4272312634;
        test_addr[2558] = 1020;
        test_data[2558] = 33'd1493206180;
        test_addr[2559] = 1021;
        test_data[2559] = 33'd349429309;
        test_addr[2560] = 1022;
        test_data[2560] = 33'd4560181166;
        test_addr[2561] = 1023;
        test_data[2561] = 33'd1545197175;
        test_addr[2562] = 0;
        test_data[2562] = 33'd1052567479;
        test_addr[2563] = 1;
        test_data[2563] = 33'd6595768149;
        test_addr[2564] = 2;
        test_data[2564] = 33'd455055946;
        test_addr[2565] = 309;
        test_data[2565] = 33'd4468640426;
        test_addr[2566] = 310;
        test_data[2566] = 33'd892285550;
        test_addr[2567] = 311;
        test_data[2567] = 33'd4809014040;
        test_addr[2568] = 312;
        test_data[2568] = 33'd1581510545;
        test_addr[2569] = 313;
        test_data[2569] = 33'd1075197784;
        test_addr[2570] = 314;
        test_data[2570] = 33'd3441385405;
        test_addr[2571] = 315;
        test_data[2571] = 33'd1538426196;
        test_addr[2572] = 316;
        test_data[2572] = 33'd2469986364;
        test_addr[2573] = 317;
        test_data[2573] = 33'd1407290752;
        test_addr[2574] = 318;
        test_data[2574] = 33'd3064576727;
        test_addr[2575] = 319;
        test_data[2575] = 33'd3903019567;
        test_addr[2576] = 320;
        test_data[2576] = 33'd8234317705;
        test_addr[2577] = 321;
        test_data[2577] = 33'd2227829365;
        test_addr[2578] = 322;
        test_data[2578] = 33'd5835407995;
        test_addr[2579] = 323;
        test_data[2579] = 33'd8171946952;
        test_addr[2580] = 324;
        test_data[2580] = 33'd7756291470;
        test_addr[2581] = 325;
        test_data[2581] = 33'd2573803079;
        test_addr[2582] = 326;
        test_data[2582] = 33'd3914629007;
        test_addr[2583] = 327;
        test_data[2583] = 33'd2931519176;
        test_addr[2584] = 328;
        test_data[2584] = 33'd2378604963;
        test_addr[2585] = 329;
        test_data[2585] = 33'd3283575319;
        test_addr[2586] = 811;
        test_data[2586] = 33'd500276442;
        test_addr[2587] = 812;
        test_data[2587] = 33'd2198066108;
        test_addr[2588] = 813;
        test_data[2588] = 33'd1567399322;
        test_addr[2589] = 814;
        test_data[2589] = 33'd2725263772;
        test_addr[2590] = 815;
        test_data[2590] = 33'd1840551582;
        test_addr[2591] = 816;
        test_data[2591] = 33'd2266625000;
        test_addr[2592] = 817;
        test_data[2592] = 33'd2256146945;
        test_addr[2593] = 818;
        test_data[2593] = 33'd4127540968;
        test_addr[2594] = 819;
        test_data[2594] = 33'd3076100910;
        test_addr[2595] = 820;
        test_data[2595] = 33'd4541216847;
        test_addr[2596] = 821;
        test_data[2596] = 33'd2641923197;
        test_addr[2597] = 822;
        test_data[2597] = 33'd1320572974;
        test_addr[2598] = 330;
        test_data[2598] = 33'd8332610434;
        test_addr[2599] = 331;
        test_data[2599] = 33'd4429917652;
        test_addr[2600] = 332;
        test_data[2600] = 33'd7687666706;
        test_addr[2601] = 333;
        test_data[2601] = 33'd2944611355;
        test_addr[2602] = 334;
        test_data[2602] = 33'd2841628197;
        test_addr[2603] = 335;
        test_data[2603] = 33'd98705679;
        test_addr[2604] = 336;
        test_data[2604] = 33'd745322449;
        test_addr[2605] = 337;
        test_data[2605] = 33'd4218420959;
        test_addr[2606] = 197;
        test_data[2606] = 33'd3233146207;
        test_addr[2607] = 198;
        test_data[2607] = 33'd6776761698;
        test_addr[2608] = 199;
        test_data[2608] = 33'd2854665516;
        test_addr[2609] = 200;
        test_data[2609] = 33'd178768342;
        test_addr[2610] = 201;
        test_data[2610] = 33'd3380527101;
        test_addr[2611] = 202;
        test_data[2611] = 33'd6646333835;
        test_addr[2612] = 203;
        test_data[2612] = 33'd2130719600;
        test_addr[2613] = 204;
        test_data[2613] = 33'd5817952334;
        test_addr[2614] = 338;
        test_data[2614] = 33'd2832891657;
        test_addr[2615] = 339;
        test_data[2615] = 33'd3237287086;
        test_addr[2616] = 340;
        test_data[2616] = 33'd2309224711;
        test_addr[2617] = 341;
        test_data[2617] = 33'd7223820858;
        test_addr[2618] = 342;
        test_data[2618] = 33'd3867550255;
        test_addr[2619] = 343;
        test_data[2619] = 33'd2642501263;
        test_addr[2620] = 468;
        test_data[2620] = 33'd4605482898;
        test_addr[2621] = 469;
        test_data[2621] = 33'd4275884649;
        test_addr[2622] = 344;
        test_data[2622] = 33'd100362266;
        test_addr[2623] = 345;
        test_data[2623] = 33'd84750818;
        test_addr[2624] = 346;
        test_data[2624] = 33'd6768287263;
        test_addr[2625] = 615;
        test_data[2625] = 33'd605372899;
        test_addr[2626] = 616;
        test_data[2626] = 33'd1345991342;
        test_addr[2627] = 347;
        test_data[2627] = 33'd6058926612;
        test_addr[2628] = 348;
        test_data[2628] = 33'd7705912888;
        test_addr[2629] = 349;
        test_data[2629] = 33'd2089693596;
        test_addr[2630] = 350;
        test_data[2630] = 33'd6705255373;
        test_addr[2631] = 351;
        test_data[2631] = 33'd4473351698;
        test_addr[2632] = 352;
        test_data[2632] = 33'd3385339541;
        test_addr[2633] = 353;
        test_data[2633] = 33'd2497359255;
        test_addr[2634] = 211;
        test_data[2634] = 33'd1230764576;
        test_addr[2635] = 354;
        test_data[2635] = 33'd4104199402;
        test_addr[2636] = 355;
        test_data[2636] = 33'd1103758275;
        test_addr[2637] = 356;
        test_data[2637] = 33'd328648182;
        test_addr[2638] = 357;
        test_data[2638] = 33'd6158270689;
        test_addr[2639] = 652;
        test_data[2639] = 33'd891912601;
        test_addr[2640] = 653;
        test_data[2640] = 33'd7978548142;
        test_addr[2641] = 654;
        test_data[2641] = 33'd7684777898;
        test_addr[2642] = 655;
        test_data[2642] = 33'd6804724310;
        test_addr[2643] = 656;
        test_data[2643] = 33'd756043176;
        test_addr[2644] = 657;
        test_data[2644] = 33'd668982047;
        test_addr[2645] = 658;
        test_data[2645] = 33'd2565372091;
        test_addr[2646] = 659;
        test_data[2646] = 33'd6970367893;
        test_addr[2647] = 660;
        test_data[2647] = 33'd7004734946;
        test_addr[2648] = 661;
        test_data[2648] = 33'd408333930;
        test_addr[2649] = 662;
        test_data[2649] = 33'd3582659021;
        test_addr[2650] = 663;
        test_data[2650] = 33'd1473735246;
        test_addr[2651] = 664;
        test_data[2651] = 33'd5670651089;
        test_addr[2652] = 665;
        test_data[2652] = 33'd1768918310;
        test_addr[2653] = 666;
        test_data[2653] = 33'd5304418194;
        test_addr[2654] = 667;
        test_data[2654] = 33'd2879010504;
        test_addr[2655] = 668;
        test_data[2655] = 33'd3382879701;
        test_addr[2656] = 669;
        test_data[2656] = 33'd3165934849;
        test_addr[2657] = 670;
        test_data[2657] = 33'd4826551882;
        test_addr[2658] = 358;
        test_data[2658] = 33'd2281669903;
        test_addr[2659] = 359;
        test_data[2659] = 33'd5777571266;
        test_addr[2660] = 360;
        test_data[2660] = 33'd1685941148;
        test_addr[2661] = 361;
        test_data[2661] = 33'd1230104128;
        test_addr[2662] = 362;
        test_data[2662] = 33'd2761902832;
        test_addr[2663] = 363;
        test_data[2663] = 33'd803716268;
        test_addr[2664] = 364;
        test_data[2664] = 33'd3270560608;
        test_addr[2665] = 365;
        test_data[2665] = 33'd6798862133;
        test_addr[2666] = 366;
        test_data[2666] = 33'd5947508543;
        test_addr[2667] = 367;
        test_data[2667] = 33'd3378755930;
        test_addr[2668] = 368;
        test_data[2668] = 33'd4912733960;
        test_addr[2669] = 369;
        test_data[2669] = 33'd2921962052;
        test_addr[2670] = 370;
        test_data[2670] = 33'd4390058828;
        test_addr[2671] = 371;
        test_data[2671] = 33'd338135865;
        test_addr[2672] = 372;
        test_data[2672] = 33'd605321337;
        test_addr[2673] = 373;
        test_data[2673] = 33'd1524839362;
        test_addr[2674] = 859;
        test_data[2674] = 33'd61833049;
        test_addr[2675] = 860;
        test_data[2675] = 33'd7160689490;
        test_addr[2676] = 861;
        test_data[2676] = 33'd4818724234;
        test_addr[2677] = 862;
        test_data[2677] = 33'd5468858884;
        test_addr[2678] = 863;
        test_data[2678] = 33'd1939476593;
        test_addr[2679] = 864;
        test_data[2679] = 33'd7875939957;
        test_addr[2680] = 374;
        test_data[2680] = 33'd3597032391;
        test_addr[2681] = 375;
        test_data[2681] = 33'd86563587;
        test_addr[2682] = 376;
        test_data[2682] = 33'd2007598323;
        test_addr[2683] = 377;
        test_data[2683] = 33'd7277834310;
        test_addr[2684] = 378;
        test_data[2684] = 33'd1683535556;
        test_addr[2685] = 724;
        test_data[2685] = 33'd3065873517;
        test_addr[2686] = 725;
        test_data[2686] = 33'd4231348663;
        test_addr[2687] = 726;
        test_data[2687] = 33'd4297080980;
        test_addr[2688] = 727;
        test_data[2688] = 33'd7262561752;
        test_addr[2689] = 728;
        test_data[2689] = 33'd3542905408;
        test_addr[2690] = 729;
        test_data[2690] = 33'd1951530555;
        test_addr[2691] = 730;
        test_data[2691] = 33'd1460298641;
        test_addr[2692] = 731;
        test_data[2692] = 33'd973228329;
        test_addr[2693] = 732;
        test_data[2693] = 33'd7919742694;
        test_addr[2694] = 733;
        test_data[2694] = 33'd2291561714;
        test_addr[2695] = 734;
        test_data[2695] = 33'd6044284591;
        test_addr[2696] = 735;
        test_data[2696] = 33'd894928856;
        test_addr[2697] = 736;
        test_data[2697] = 33'd5906561941;
        test_addr[2698] = 379;
        test_data[2698] = 33'd2072366047;
        test_addr[2699] = 227;
        test_data[2699] = 33'd6767044533;
        test_addr[2700] = 228;
        test_data[2700] = 33'd1793161912;
        test_addr[2701] = 229;
        test_data[2701] = 33'd1524904068;
        test_addr[2702] = 230;
        test_data[2702] = 33'd1629741321;
        test_addr[2703] = 231;
        test_data[2703] = 33'd6669555233;
        test_addr[2704] = 232;
        test_data[2704] = 33'd274384184;
        test_addr[2705] = 233;
        test_data[2705] = 33'd312253816;
        test_addr[2706] = 234;
        test_data[2706] = 33'd4056501288;
        test_addr[2707] = 235;
        test_data[2707] = 33'd5152104255;
        test_addr[2708] = 236;
        test_data[2708] = 33'd2037725383;
        test_addr[2709] = 237;
        test_data[2709] = 33'd1838823857;
        test_addr[2710] = 238;
        test_data[2710] = 33'd3263906087;
        test_addr[2711] = 239;
        test_data[2711] = 33'd935814712;
        test_addr[2712] = 240;
        test_data[2712] = 33'd1543222631;
        test_addr[2713] = 241;
        test_data[2713] = 33'd3949767492;
        test_addr[2714] = 380;
        test_data[2714] = 33'd4349868449;
        test_addr[2715] = 381;
        test_data[2715] = 33'd1148986808;
        test_addr[2716] = 382;
        test_data[2716] = 33'd4817776623;
        test_addr[2717] = 383;
        test_data[2717] = 33'd51573383;
        test_addr[2718] = 384;
        test_data[2718] = 33'd1409343159;
        test_addr[2719] = 385;
        test_data[2719] = 33'd5590630983;
        test_addr[2720] = 386;
        test_data[2720] = 33'd5091387776;
        test_addr[2721] = 387;
        test_data[2721] = 33'd4976428597;
        test_addr[2722] = 388;
        test_data[2722] = 33'd222049690;
        test_addr[2723] = 325;
        test_data[2723] = 33'd8234995887;
        test_addr[2724] = 326;
        test_data[2724] = 33'd3914629007;
        test_addr[2725] = 327;
        test_data[2725] = 33'd5703386628;
        test_addr[2726] = 328;
        test_data[2726] = 33'd2378604963;
        test_addr[2727] = 329;
        test_data[2727] = 33'd3283575319;
        test_addr[2728] = 330;
        test_data[2728] = 33'd6392011536;
        test_addr[2729] = 331;
        test_data[2729] = 33'd4976018475;
        test_addr[2730] = 332;
        test_data[2730] = 33'd3392699410;
        test_addr[2731] = 333;
        test_data[2731] = 33'd2944611355;
        test_addr[2732] = 334;
        test_data[2732] = 33'd2841628197;
        test_addr[2733] = 335;
        test_data[2733] = 33'd98705679;
        test_addr[2734] = 336;
        test_data[2734] = 33'd745322449;
        test_addr[2735] = 337;
        test_data[2735] = 33'd7289977960;
        test_addr[2736] = 338;
        test_data[2736] = 33'd8083651609;
        test_addr[2737] = 339;
        test_data[2737] = 33'd3237287086;
        test_addr[2738] = 340;
        test_data[2738] = 33'd2309224711;
        test_addr[2739] = 341;
        test_data[2739] = 33'd6418123408;
        test_addr[2740] = 342;
        test_data[2740] = 33'd3867550255;
        test_addr[2741] = 343;
        test_data[2741] = 33'd2642501263;
        test_addr[2742] = 344;
        test_data[2742] = 33'd5552826033;
        test_addr[2743] = 345;
        test_data[2743] = 33'd6807917029;
        test_addr[2744] = 346;
        test_data[2744] = 33'd2473319967;
        test_addr[2745] = 347;
        test_data[2745] = 33'd1763959316;
        test_addr[2746] = 348;
        test_data[2746] = 33'd3410945592;
        test_addr[2747] = 349;
        test_data[2747] = 33'd2089693596;
        test_addr[2748] = 350;
        test_data[2748] = 33'd2410288077;
        test_addr[2749] = 351;
        test_data[2749] = 33'd178384402;
        test_addr[2750] = 352;
        test_data[2750] = 33'd3385339541;
        test_addr[2751] = 353;
        test_data[2751] = 33'd2497359255;
        test_addr[2752] = 354;
        test_data[2752] = 33'd7246375191;
        test_addr[2753] = 355;
        test_data[2753] = 33'd1103758275;
        test_addr[2754] = 389;
        test_data[2754] = 33'd4280400511;
        test_addr[2755] = 390;
        test_data[2755] = 33'd4980712302;
        test_addr[2756] = 391;
        test_data[2756] = 33'd22882165;
        test_addr[2757] = 392;
        test_data[2757] = 33'd2454339683;
        test_addr[2758] = 931;
        test_data[2758] = 33'd7928129;
        test_addr[2759] = 932;
        test_data[2759] = 33'd1498951355;
        test_addr[2760] = 933;
        test_data[2760] = 33'd5702913498;
        test_addr[2761] = 934;
        test_data[2761] = 33'd5175624083;
        test_addr[2762] = 935;
        test_data[2762] = 33'd3119130326;
        test_addr[2763] = 936;
        test_data[2763] = 33'd4710482889;
        test_addr[2764] = 937;
        test_data[2764] = 33'd7885826526;
        test_addr[2765] = 393;
        test_data[2765] = 33'd3236922202;
        test_addr[2766] = 394;
        test_data[2766] = 33'd5452117273;
        test_addr[2767] = 395;
        test_data[2767] = 33'd101142806;
        test_addr[2768] = 396;
        test_data[2768] = 33'd3707484179;
        test_addr[2769] = 397;
        test_data[2769] = 33'd6801216116;
        test_addr[2770] = 398;
        test_data[2770] = 33'd3583158237;
        test_addr[2771] = 399;
        test_data[2771] = 33'd6742062650;
        test_addr[2772] = 400;
        test_data[2772] = 33'd4549000436;
        test_addr[2773] = 401;
        test_data[2773] = 33'd7103521096;
        test_addr[2774] = 402;
        test_data[2774] = 33'd1240298673;
        test_addr[2775] = 403;
        test_data[2775] = 33'd7346723591;
        test_addr[2776] = 404;
        test_data[2776] = 33'd2974441075;
        test_addr[2777] = 405;
        test_data[2777] = 33'd5550819530;
        test_addr[2778] = 406;
        test_data[2778] = 33'd5430851424;
        test_addr[2779] = 407;
        test_data[2779] = 33'd4772195850;
        test_addr[2780] = 408;
        test_data[2780] = 33'd2708666325;
        test_addr[2781] = 43;
        test_data[2781] = 33'd2262236211;
        test_addr[2782] = 44;
        test_data[2782] = 33'd1578693673;
        test_addr[2783] = 45;
        test_data[2783] = 33'd3465150654;
        test_addr[2784] = 46;
        test_data[2784] = 33'd3718565962;
        test_addr[2785] = 47;
        test_data[2785] = 33'd7903934043;
        test_addr[2786] = 409;
        test_data[2786] = 33'd664332654;
        test_addr[2787] = 410;
        test_data[2787] = 33'd2554823396;
        test_addr[2788] = 411;
        test_data[2788] = 33'd7395462392;
        test_addr[2789] = 412;
        test_data[2789] = 33'd1136766050;
        test_addr[2790] = 413;
        test_data[2790] = 33'd42785687;
        test_addr[2791] = 414;
        test_data[2791] = 33'd650430649;
        test_addr[2792] = 415;
        test_data[2792] = 33'd7196900617;
        test_addr[2793] = 416;
        test_data[2793] = 33'd6253627735;
        test_addr[2794] = 417;
        test_data[2794] = 33'd3609631975;
        test_addr[2795] = 38;
        test_data[2795] = 33'd982384382;
        test_addr[2796] = 39;
        test_data[2796] = 33'd1162677645;
        test_addr[2797] = 40;
        test_data[2797] = 33'd334310572;
        test_addr[2798] = 41;
        test_data[2798] = 33'd897063482;
        test_addr[2799] = 42;
        test_data[2799] = 33'd7546933915;
        test_addr[2800] = 43;
        test_data[2800] = 33'd6218261399;
        test_addr[2801] = 44;
        test_data[2801] = 33'd1578693673;
        test_addr[2802] = 45;
        test_data[2802] = 33'd8046824005;
        test_addr[2803] = 46;
        test_data[2803] = 33'd3718565962;
        test_addr[2804] = 47;
        test_data[2804] = 33'd5999281312;
        test_addr[2805] = 48;
        test_data[2805] = 33'd8028059791;
        test_addr[2806] = 49;
        test_data[2806] = 33'd453190497;
        test_addr[2807] = 50;
        test_data[2807] = 33'd304764150;
        test_addr[2808] = 51;
        test_data[2808] = 33'd2861275312;
        test_addr[2809] = 52;
        test_data[2809] = 33'd2084213537;
        test_addr[2810] = 53;
        test_data[2810] = 33'd5658971079;
        test_addr[2811] = 54;
        test_data[2811] = 33'd255843487;
        test_addr[2812] = 418;
        test_data[2812] = 33'd440038134;
        test_addr[2813] = 419;
        test_data[2813] = 33'd6718911545;
        test_addr[2814] = 420;
        test_data[2814] = 33'd7335937971;
        test_addr[2815] = 421;
        test_data[2815] = 33'd749396176;
        test_addr[2816] = 422;
        test_data[2816] = 33'd4129404128;
        test_addr[2817] = 423;
        test_data[2817] = 33'd6411449459;
        test_addr[2818] = 428;
        test_data[2818] = 33'd3112127436;
        test_addr[2819] = 429;
        test_data[2819] = 33'd496696578;
        test_addr[2820] = 430;
        test_data[2820] = 33'd3912201120;
        test_addr[2821] = 431;
        test_data[2821] = 33'd2084255774;
        test_addr[2822] = 432;
        test_data[2822] = 33'd807161466;
        test_addr[2823] = 433;
        test_data[2823] = 33'd363795349;
        test_addr[2824] = 434;
        test_data[2824] = 33'd2998754042;
        test_addr[2825] = 435;
        test_data[2825] = 33'd6791735478;
        test_addr[2826] = 436;
        test_data[2826] = 33'd4273322909;
        test_addr[2827] = 437;
        test_data[2827] = 33'd1332405155;
        test_addr[2828] = 438;
        test_data[2828] = 33'd2165787536;
        test_addr[2829] = 439;
        test_data[2829] = 33'd6840001730;
        test_addr[2830] = 440;
        test_data[2830] = 33'd3037982191;
        test_addr[2831] = 441;
        test_data[2831] = 33'd7546066905;
        test_addr[2832] = 442;
        test_data[2832] = 33'd4170323346;
        test_addr[2833] = 443;
        test_data[2833] = 33'd1076063113;
        test_addr[2834] = 444;
        test_data[2834] = 33'd4084632541;
        test_addr[2835] = 445;
        test_data[2835] = 33'd1727324708;
        test_addr[2836] = 446;
        test_data[2836] = 33'd2468389652;
        test_addr[2837] = 447;
        test_data[2837] = 33'd3376647238;
        test_addr[2838] = 448;
        test_data[2838] = 33'd7977205554;
        test_addr[2839] = 424;
        test_data[2839] = 33'd4259167484;
        test_addr[2840] = 425;
        test_data[2840] = 33'd3432594820;
        test_addr[2841] = 426;
        test_data[2841] = 33'd6910994609;
        test_addr[2842] = 427;
        test_data[2842] = 33'd3990194643;
        test_addr[2843] = 428;
        test_data[2843] = 33'd5595175681;
        test_addr[2844] = 429;
        test_data[2844] = 33'd496696578;
        test_addr[2845] = 430;
        test_data[2845] = 33'd3912201120;
        test_addr[2846] = 431;
        test_data[2846] = 33'd2084255774;
        test_addr[2847] = 432;
        test_data[2847] = 33'd807161466;
        test_addr[2848] = 433;
        test_data[2848] = 33'd8408494181;
        test_addr[2849] = 434;
        test_data[2849] = 33'd2998754042;
        test_addr[2850] = 435;
        test_data[2850] = 33'd2496768182;
        test_addr[2851] = 436;
        test_data[2851] = 33'd7773873709;
        test_addr[2852] = 437;
        test_data[2852] = 33'd1332405155;
        test_addr[2853] = 438;
        test_data[2853] = 33'd6793367620;
        test_addr[2854] = 439;
        test_data[2854] = 33'd2545034434;
        test_addr[2855] = 440;
        test_data[2855] = 33'd3037982191;
        test_addr[2856] = 441;
        test_data[2856] = 33'd3251099609;
        test_addr[2857] = 442;
        test_data[2857] = 33'd4170323346;
        test_addr[2858] = 443;
        test_data[2858] = 33'd6560361925;
        test_addr[2859] = 444;
        test_data[2859] = 33'd4084632541;
        test_addr[2860] = 445;
        test_data[2860] = 33'd1727324708;
        test_addr[2861] = 446;
        test_data[2861] = 33'd2468389652;
        test_addr[2862] = 447;
        test_data[2862] = 33'd3376647238;
        test_addr[2863] = 448;
        test_data[2863] = 33'd3682238258;
        test_addr[2864] = 449;
        test_data[2864] = 33'd2908833870;
        test_addr[2865] = 450;
        test_data[2865] = 33'd2162667854;
        test_addr[2866] = 451;
        test_data[2866] = 33'd3487811640;
        test_addr[2867] = 452;
        test_data[2867] = 33'd548840626;
        test_addr[2868] = 453;
        test_data[2868] = 33'd7583003951;
        test_addr[2869] = 454;
        test_data[2869] = 33'd1295592959;
        test_addr[2870] = 455;
        test_data[2870] = 33'd2580577157;
        test_addr[2871] = 456;
        test_data[2871] = 33'd5050570264;
        test_addr[2872] = 457;
        test_data[2872] = 33'd6684942309;
        test_addr[2873] = 458;
        test_data[2873] = 33'd5160448221;
        test_addr[2874] = 459;
        test_data[2874] = 33'd6087096786;
        test_addr[2875] = 460;
        test_data[2875] = 33'd2220856156;
        test_addr[2876] = 461;
        test_data[2876] = 33'd3428994727;
        test_addr[2877] = 462;
        test_data[2877] = 33'd151052727;
        test_addr[2878] = 463;
        test_data[2878] = 33'd1720502167;
        test_addr[2879] = 464;
        test_data[2879] = 33'd1825193099;
        test_addr[2880] = 465;
        test_data[2880] = 33'd3508624685;
        test_addr[2881] = 466;
        test_data[2881] = 33'd1761019531;
        test_addr[2882] = 467;
        test_data[2882] = 33'd1066574642;
        test_addr[2883] = 468;
        test_data[2883] = 33'd310515602;
        test_addr[2884] = 469;
        test_data[2884] = 33'd4275884649;
        test_addr[2885] = 470;
        test_data[2885] = 33'd8373215536;
        test_addr[2886] = 471;
        test_data[2886] = 33'd996654737;
        test_addr[2887] = 472;
        test_data[2887] = 33'd173483137;
        test_addr[2888] = 797;
        test_data[2888] = 33'd3100043597;
        test_addr[2889] = 798;
        test_data[2889] = 33'd3715808831;
        test_addr[2890] = 799;
        test_data[2890] = 33'd4174440399;
        test_addr[2891] = 800;
        test_data[2891] = 33'd356101764;
        test_addr[2892] = 801;
        test_data[2892] = 33'd4030133163;
        test_addr[2893] = 802;
        test_data[2893] = 33'd6558952631;
        test_addr[2894] = 803;
        test_data[2894] = 33'd3130885866;
        test_addr[2895] = 804;
        test_data[2895] = 33'd8448614737;
        test_addr[2896] = 805;
        test_data[2896] = 33'd4670308951;
        test_addr[2897] = 806;
        test_data[2897] = 33'd2394794120;
        test_addr[2898] = 473;
        test_data[2898] = 33'd6782211258;
        test_addr[2899] = 474;
        test_data[2899] = 33'd3821064159;
        test_addr[2900] = 475;
        test_data[2900] = 33'd3328634438;
        test_addr[2901] = 476;
        test_data[2901] = 33'd7891126102;
        test_addr[2902] = 477;
        test_data[2902] = 33'd7348033864;
        test_addr[2903] = 478;
        test_data[2903] = 33'd5776234055;
        test_addr[2904] = 479;
        test_data[2904] = 33'd2293417793;
        test_addr[2905] = 480;
        test_data[2905] = 33'd799026300;
        test_addr[2906] = 481;
        test_data[2906] = 33'd3611509395;
        test_addr[2907] = 971;
        test_data[2907] = 33'd7841993419;
        test_addr[2908] = 972;
        test_data[2908] = 33'd1407407298;
        test_addr[2909] = 482;
        test_data[2909] = 33'd6356614554;
        test_addr[2910] = 483;
        test_data[2910] = 33'd2772842294;
        test_addr[2911] = 586;
        test_data[2911] = 33'd3351735354;
        test_addr[2912] = 587;
        test_data[2912] = 33'd291280601;
        test_addr[2913] = 588;
        test_data[2913] = 33'd4621878581;
        test_addr[2914] = 484;
        test_data[2914] = 33'd4037018018;
        test_addr[2915] = 485;
        test_data[2915] = 33'd453359906;
        test_addr[2916] = 486;
        test_data[2916] = 33'd6610140484;
        test_addr[2917] = 487;
        test_data[2917] = 33'd3658540064;
        test_addr[2918] = 488;
        test_data[2918] = 33'd2552432527;
        test_addr[2919] = 489;
        test_data[2919] = 33'd1327010194;
        test_addr[2920] = 1001;
        test_data[2920] = 33'd2748983834;
        test_addr[2921] = 1002;
        test_data[2921] = 33'd1328575902;
        test_addr[2922] = 1003;
        test_data[2922] = 33'd7529868376;
        test_addr[2923] = 1004;
        test_data[2923] = 33'd784496299;
        test_addr[2924] = 1005;
        test_data[2924] = 33'd3407483378;
        test_addr[2925] = 1006;
        test_data[2925] = 33'd1958914203;
        test_addr[2926] = 1007;
        test_data[2926] = 33'd5919413050;
        test_addr[2927] = 1008;
        test_data[2927] = 33'd457320104;
        test_addr[2928] = 1009;
        test_data[2928] = 33'd3497266080;
        test_addr[2929] = 1010;
        test_data[2929] = 33'd3905914762;
        test_addr[2930] = 1011;
        test_data[2930] = 33'd2784490477;
        test_addr[2931] = 1012;
        test_data[2931] = 33'd7817989407;
        test_addr[2932] = 1013;
        test_data[2932] = 33'd6427759724;
        test_addr[2933] = 490;
        test_data[2933] = 33'd1847146603;
        test_addr[2934] = 491;
        test_data[2934] = 33'd7281999275;
        test_addr[2935] = 492;
        test_data[2935] = 33'd5860388549;
        test_addr[2936] = 493;
        test_data[2936] = 33'd909000303;
        test_addr[2937] = 494;
        test_data[2937] = 33'd5183494673;
        test_addr[2938] = 495;
        test_data[2938] = 33'd3025805301;
        test_addr[2939] = 496;
        test_data[2939] = 33'd3017411151;
        test_addr[2940] = 497;
        test_data[2940] = 33'd6298676298;
        test_addr[2941] = 498;
        test_data[2941] = 33'd4345254171;
        test_addr[2942] = 499;
        test_data[2942] = 33'd1806570311;
        test_addr[2943] = 500;
        test_data[2943] = 33'd1186374242;
        test_addr[2944] = 501;
        test_data[2944] = 33'd2724914268;
        test_addr[2945] = 502;
        test_data[2945] = 33'd6012534491;
        test_addr[2946] = 503;
        test_data[2946] = 33'd4493817892;
        test_addr[2947] = 504;
        test_data[2947] = 33'd1574083226;
        test_addr[2948] = 505;
        test_data[2948] = 33'd3026237748;
        test_addr[2949] = 506;
        test_data[2949] = 33'd307644181;
        test_addr[2950] = 507;
        test_data[2950] = 33'd2717188915;
        test_addr[2951] = 508;
        test_data[2951] = 33'd7250565982;
        test_addr[2952] = 509;
        test_data[2952] = 33'd282828349;
        test_addr[2953] = 220;
        test_data[2953] = 33'd7292249776;
        test_addr[2954] = 221;
        test_data[2954] = 33'd2513170581;
        test_addr[2955] = 222;
        test_data[2955] = 33'd3954542123;
        test_addr[2956] = 223;
        test_data[2956] = 33'd1645865683;
        test_addr[2957] = 224;
        test_data[2957] = 33'd11908938;
        test_addr[2958] = 225;
        test_data[2958] = 33'd8129806786;
        test_addr[2959] = 226;
        test_data[2959] = 33'd4073331549;
        test_addr[2960] = 227;
        test_data[2960] = 33'd2472077237;
        test_addr[2961] = 228;
        test_data[2961] = 33'd1793161912;
        test_addr[2962] = 229;
        test_data[2962] = 33'd1524904068;
        test_addr[2963] = 230;
        test_data[2963] = 33'd1629741321;
        test_addr[2964] = 231;
        test_data[2964] = 33'd4626792729;
        test_addr[2965] = 232;
        test_data[2965] = 33'd274384184;
        test_addr[2966] = 233;
        test_data[2966] = 33'd7056180896;
        test_addr[2967] = 234;
        test_data[2967] = 33'd8372843144;
        test_addr[2968] = 235;
        test_data[2968] = 33'd857136959;
        test_addr[2969] = 236;
        test_data[2969] = 33'd6281745466;
        test_addr[2970] = 237;
        test_data[2970] = 33'd1838823857;
        test_addr[2971] = 238;
        test_data[2971] = 33'd3263906087;
        test_addr[2972] = 239;
        test_data[2972] = 33'd4635109738;
        test_addr[2973] = 240;
        test_data[2973] = 33'd6502304274;
        test_addr[2974] = 241;
        test_data[2974] = 33'd3949767492;
        test_addr[2975] = 242;
        test_data[2975] = 33'd136386603;
        test_addr[2976] = 510;
        test_data[2976] = 33'd4584807539;
        test_addr[2977] = 511;
        test_data[2977] = 33'd6838572878;
        test_addr[2978] = 206;
        test_data[2978] = 33'd1500141252;
        test_addr[2979] = 207;
        test_data[2979] = 33'd6510060590;
        test_addr[2980] = 208;
        test_data[2980] = 33'd5054016943;
        test_addr[2981] = 209;
        test_data[2981] = 33'd4188964105;
        test_addr[2982] = 512;
        test_data[2982] = 33'd1811787911;
        test_addr[2983] = 513;
        test_data[2983] = 33'd6492642645;
        test_addr[2984] = 514;
        test_data[2984] = 33'd2760410661;
        test_addr[2985] = 515;
        test_data[2985] = 33'd3342319872;
        test_addr[2986] = 880;
        test_data[2986] = 33'd830185165;
        test_addr[2987] = 881;
        test_data[2987] = 33'd1506016935;
        test_addr[2988] = 882;
        test_data[2988] = 33'd3835130572;
        test_addr[2989] = 883;
        test_data[2989] = 33'd3004317571;
        test_addr[2990] = 884;
        test_data[2990] = 33'd422576570;
        test_addr[2991] = 885;
        test_data[2991] = 33'd2842593496;
        test_addr[2992] = 886;
        test_data[2992] = 33'd377684310;
        test_addr[2993] = 887;
        test_data[2993] = 33'd3092087050;
        test_addr[2994] = 888;
        test_data[2994] = 33'd309666434;
        test_addr[2995] = 889;
        test_data[2995] = 33'd2093999100;
        test_addr[2996] = 890;
        test_data[2996] = 33'd1874897802;
        test_addr[2997] = 891;
        test_data[2997] = 33'd4360217858;
        test_addr[2998] = 516;
        test_data[2998] = 33'd6958703378;
        test_addr[2999] = 517;
        test_data[2999] = 33'd5380495514;

    end
endmodule
